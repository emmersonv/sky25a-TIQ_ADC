magic
tech sky130A
timestamp 1754266322
<< nwell >>
rect 131 461 153 479
rect 262 461 284 479
rect 113 361 171 461
rect 244 361 302 461
rect 131 203 153 361
rect 262 203 284 361
<< nsubdiff >>
rect 113 361 171 461
rect 244 361 302 461
<< locali >>
rect 0 195 8 202
rect 385 194 393 201
<< metal1 >>
rect 185 446 202 454
rect 186 8 203 16
use inverter_p1_n0o42  inverter_p1_n0o42_0
timestamp 1754263527
transform 1 0 40 0 1 114
box -40 -114 91 365
use inverter_p1_n0o42  inverter_p1_n0o42_1
timestamp 1754263527
transform 1 0 171 0 1 114
box -40 -114 91 365
use inverter_p1_n0o42  inverter_p1_n0o42_2
timestamp 1754263527
transform 1 0 302 0 1 114
box -40 -114 91 365
<< labels >>
rlabel locali 0 195 8 202 7 in
port 1 w
rlabel locali 385 194 393 201 3 out
port 2 e
rlabel metal1 186 8 203 16 5 VGND
port 3 s
rlabel metal1 185 446 202 454 1 VDPWR
port 4 n
<< end >>
