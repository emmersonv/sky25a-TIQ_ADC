magic
tech sky130A
magscale 1 2
timestamp 1756008383
<< error_s >>
rect 4900 4300 5100 4458
rect 5136 4300 5268 4468
rect 4900 4264 5268 4300
rect 5100 4240 5268 4264
rect 4900 4204 5268 4240
rect 4900 4168 5100 4204
<< locali >>
rect 208 6319 274 6336
rect 208 6285 224 6319
rect 258 6285 274 6319
rect 208 6268 274 6285
rect 208 5333 274 5348
rect 208 5299 224 5333
rect 258 5299 274 5333
rect 208 5280 274 5299
rect 208 4349 274 4366
rect 208 4315 224 4349
rect 258 4315 274 4349
rect 208 4298 274 4315
rect 208 3365 274 3382
rect 208 3331 224 3365
rect 258 3331 274 3365
rect 208 3314 274 3331
rect 208 2381 274 2398
rect 208 2347 224 2381
rect 258 2347 274 2381
rect 208 2330 274 2347
rect 208 1395 274 1412
rect 208 1361 224 1395
rect 258 1361 274 1395
rect 208 1344 274 1361
rect 208 411 274 428
rect 208 377 224 411
rect 258 377 274 411
rect 208 360 274 377
<< viali >>
rect 224 6285 258 6319
rect 224 5299 258 5333
rect 224 4315 258 4349
rect 224 3331 258 3365
rect 224 2347 258 2381
rect 224 1361 258 1395
rect 224 377 258 411
<< metal1 >>
rect -130 6814 5082 6820
rect -3860 6805 5082 6814
rect -3860 6753 -3849 6805
rect -3797 6753 -3769 6805
rect -3717 6753 -3689 6805
rect -3637 6753 -3609 6805
rect -3557 6753 5082 6805
rect -3860 6725 5082 6753
rect -3860 6673 -3849 6725
rect -3797 6673 -3769 6725
rect -3717 6673 -3689 6725
rect -3637 6673 -3609 6725
rect -3557 6673 5082 6725
rect -3860 6640 5082 6673
rect -130 6638 5082 6640
rect 208 6329 274 6336
rect 208 6277 215 6329
rect 267 6277 274 6329
rect 208 6268 274 6277
rect 208 5341 274 5348
rect 208 5289 215 5341
rect 267 5289 274 5341
rect 208 5280 274 5289
rect 208 4359 274 4366
rect 208 4307 215 4359
rect 267 4307 274 4359
rect 208 4298 274 4307
rect 208 3375 274 3382
rect 208 3323 215 3375
rect 267 3323 274 3375
rect 208 3314 274 3323
rect 208 2391 274 2398
rect 208 2339 215 2391
rect 267 2339 274 2391
rect 208 2330 274 2339
rect 208 1405 274 1412
rect 208 1353 215 1405
rect 267 1353 274 1405
rect 208 1344 274 1353
rect 208 421 274 428
rect 208 369 215 421
rect 267 369 274 421
rect 208 360 274 369
rect -3200 155 1324 184
rect -3200 103 -3187 155
rect -3135 103 -3107 155
rect -3055 103 -3027 155
rect -2975 103 -2947 155
rect -2895 103 1324 155
rect -3200 75 1324 103
rect -3200 23 -3187 75
rect -3135 23 -3107 75
rect -3055 23 -3027 75
rect -2975 23 -2947 75
rect -2895 23 1324 75
rect -3200 16 1324 23
<< via1 >>
rect -3849 6753 -3797 6805
rect -3769 6753 -3717 6805
rect -3689 6753 -3637 6805
rect -3609 6753 -3557 6805
rect -3849 6673 -3797 6725
rect -3769 6673 -3717 6725
rect -3689 6673 -3637 6725
rect -3609 6673 -3557 6725
rect 215 6319 267 6329
rect 215 6285 224 6319
rect 224 6285 258 6319
rect 258 6285 267 6319
rect 215 6277 267 6285
rect 215 5333 267 5341
rect 215 5299 224 5333
rect 224 5299 258 5333
rect 258 5299 267 5333
rect 215 5289 267 5299
rect 215 4349 267 4359
rect 215 4315 224 4349
rect 224 4315 258 4349
rect 258 4315 267 4349
rect 215 4307 267 4315
rect 215 3365 267 3375
rect 215 3331 224 3365
rect 224 3331 258 3365
rect 258 3331 267 3365
rect 215 3323 267 3331
rect 215 2381 267 2391
rect 215 2347 224 2381
rect 224 2347 258 2381
rect 258 2347 267 2381
rect 215 2339 267 2347
rect 215 1395 267 1405
rect 215 1361 224 1395
rect 224 1361 258 1395
rect 258 1361 267 1395
rect 215 1353 267 1361
rect 215 411 267 421
rect 215 377 224 411
rect 224 377 258 411
rect 258 377 267 411
rect 215 369 267 377
rect -3187 103 -3135 155
rect -3107 103 -3055 155
rect -3027 103 -2975 155
rect -2947 103 -2895 155
rect -3187 23 -3135 75
rect -3107 23 -3055 75
rect -3027 23 -2975 75
rect -2947 23 -2895 75
<< metal2 >>
rect -260 6818 -192 6828
rect -3860 6808 -3540 6814
rect -3860 6672 -3850 6808
rect -3554 6672 -3540 6808
rect -3860 6640 -3540 6672
rect -260 6762 -254 6818
rect -198 6762 -192 6818
rect -260 6336 -192 6762
rect -260 6329 274 6336
rect -260 6277 215 6329
rect 267 6277 274 6329
rect -260 6268 274 6277
rect -238 5732 -170 5742
rect -238 5676 -232 5732
rect -176 5676 -170 5732
rect -238 5348 -170 5676
rect -238 5341 274 5348
rect -238 5289 215 5341
rect 267 5289 274 5341
rect -238 5280 274 5289
rect -238 4644 -170 4654
rect -238 4588 -232 4644
rect -176 4588 -170 4644
rect -238 4366 -170 4588
rect -238 4359 274 4366
rect -238 4307 215 4359
rect 267 4307 274 4359
rect -238 4298 274 4307
rect -238 3558 -170 3568
rect -238 3502 -232 3558
rect -176 3502 -170 3558
rect 2862 3506 2896 3664
rect -238 3382 -170 3502
rect -238 3375 274 3382
rect -238 3323 215 3375
rect 267 3323 274 3375
rect -238 3314 274 3323
rect -238 2462 -170 2472
rect -238 2406 -232 2462
rect -176 2406 -170 2462
rect -238 2398 -170 2406
rect -238 2391 274 2398
rect -238 2339 215 2391
rect 267 2339 274 2391
rect -238 2330 274 2339
rect -238 1405 274 1412
rect -238 1384 215 1405
rect -238 1328 -232 1384
rect -176 1353 215 1384
rect 267 1353 274 1405
rect -176 1344 274 1353
rect -176 1328 -170 1344
rect -238 1314 -170 1328
rect -3818 324 -3762 1016
rect -238 421 274 428
rect -238 369 215 421
rect 267 369 274 421
rect -238 360 274 369
rect -238 298 -170 360
rect -238 242 -232 298
rect -176 242 -170 298
rect -238 232 -170 242
rect -3200 158 -2880 184
rect -3200 22 -3188 158
rect -2892 22 -2880 158
rect -3200 16 -2880 22
<< via2 >>
rect -3850 6805 -3554 6808
rect -3850 6753 -3849 6805
rect -3849 6753 -3797 6805
rect -3797 6753 -3769 6805
rect -3769 6753 -3717 6805
rect -3717 6753 -3689 6805
rect -3689 6753 -3637 6805
rect -3637 6753 -3609 6805
rect -3609 6753 -3557 6805
rect -3557 6753 -3554 6805
rect -3850 6725 -3554 6753
rect -3850 6673 -3849 6725
rect -3849 6673 -3797 6725
rect -3797 6673 -3769 6725
rect -3769 6673 -3717 6725
rect -3717 6673 -3689 6725
rect -3689 6673 -3637 6725
rect -3637 6673 -3609 6725
rect -3609 6673 -3557 6725
rect -3557 6673 -3554 6725
rect -3850 6672 -3554 6673
rect -254 6762 -198 6818
rect -232 5676 -176 5732
rect -232 4588 -176 4644
rect -232 3502 -176 3558
rect -232 2406 -176 2462
rect -232 1328 -176 1384
rect -232 242 -176 298
rect -3188 155 -2892 158
rect -3188 103 -3187 155
rect -3187 103 -3135 155
rect -3135 103 -3107 155
rect -3107 103 -3055 155
rect -3055 103 -3027 155
rect -3027 103 -2975 155
rect -2975 103 -2947 155
rect -2947 103 -2895 155
rect -2895 103 -2892 155
rect -3188 75 -2892 103
rect -3188 23 -3187 75
rect -3187 23 -3135 75
rect -3135 23 -3107 75
rect -3107 23 -3055 75
rect -3055 23 -3027 75
rect -3027 23 -2975 75
rect -2975 23 -2947 75
rect -2947 23 -2895 75
rect -2895 23 -2892 75
rect -3188 22 -2892 23
<< metal3 >>
rect -276 6818 -178 6840
rect -3860 6812 -3540 6814
rect -3860 6668 -3854 6812
rect -3550 6668 -3540 6812
rect -276 6762 -254 6818
rect -198 6762 -178 6818
rect -276 6742 -178 6762
rect -3860 6640 -3540 6668
rect -7516 5916 -7116 6036
rect -254 5732 -156 5754
rect -254 5676 -232 5732
rect -176 5676 -156 5732
rect -254 5656 -156 5676
rect -254 4644 -156 4664
rect -254 4588 -232 4644
rect -176 4588 -156 4644
rect -254 4566 -156 4588
rect -7514 3468 -7114 3588
rect -254 3558 -156 3578
rect -254 3502 -232 3558
rect -176 3502 -156 3558
rect -254 3480 -156 3502
rect -256 2462 -158 2486
rect -256 2406 -232 2462
rect -176 2406 -158 2462
rect -256 2388 -158 2406
rect -254 1384 -156 1400
rect -254 1328 -232 1384
rect -176 1328 -156 1384
rect -254 1302 -156 1328
rect -7516 1020 -7116 1140
rect -256 298 -158 316
rect -256 242 -232 298
rect -176 242 -158 298
rect -256 218 -158 242
rect -3200 162 -2880 184
rect -3200 18 -3192 162
rect -2888 18 -2880 162
rect -3200 16 -2880 18
<< via3 >>
rect -3854 6808 -3550 6812
rect -3854 6672 -3850 6808
rect -3850 6672 -3554 6808
rect -3554 6672 -3550 6808
rect -3854 6668 -3550 6672
rect -3192 158 -2888 162
rect -3192 22 -3188 158
rect -3188 22 -2892 158
rect -2892 22 -2888 158
rect -3192 18 -2888 22
<< metal4 >>
rect -3860 6812 -3540 6814
rect -3860 6668 -3854 6812
rect -3550 6668 -3540 6812
rect -3860 6500 -3540 6668
rect -3200 162 -2880 420
rect -3200 18 -3192 162
rect -2888 18 -2880 162
rect -3200 16 -2880 18
use boosted_tiq_adc_7  boosted_tiq_adc_7_0
timestamp 1756008383
transform 1 0 260 0 1 0
box -260 -26 5008 6864
use encoder  encoder_0
timestamp 1756008383
transform 1 0 -7516 0 1 -76
box 0 0 7471 6928
<< labels >>
rlabel metal1 s -548 16 -380 184 4 VGND
port 1 nsew
rlabel metal1 s -658 6640 -494 6814 4 VDPWR
port 2 nsew
rlabel metal2 s 2862 3506 2896 3664 4 Vin
port 3 nsew
rlabel metal3 s -7516 1020 -7116 1140 4 o0
port 4 nsew
rlabel metal3 s -7514 3468 -7114 3588 4 o1
port 5 nsew
rlabel metal3 s -7516 5916 -7116 6036 4 o2
port 6 nsew
<< end >>
