magic
tech sky130A
magscale 1 2
timestamp 1755919380
<< error_s >>
rect -36 3346 590 3396
rect 0 3324 554 3346
rect 0 3310 36 3324
rect 518 3310 554 3324
rect 626 3258 734 3366
rect 0 3196 36 3210
rect 518 3196 554 3210
rect 0 3174 554 3196
rect -36 3160 590 3174
rect -36 3124 172 3160
rect 206 3124 590 3160
rect 206 1654 340 3124
<< nwell >>
rect 0 3346 554 3360
rect -36 3174 590 3346
rect 0 3160 554 3174
rect 172 1646 206 3160
rect -36 1130 590 1646
<< psubdiff >>
rect 0 -432 590 -400
rect 0 -468 76 -432
rect 112 -468 168 -432
rect 204 -468 260 -432
rect 296 -468 352 -432
rect 388 -468 444 -432
rect 480 -468 536 -432
rect 572 -468 590 -432
rect 0 -524 590 -468
rect 0 -560 76 -524
rect 112 -560 168 -524
rect 204 -560 260 -524
rect 296 -560 352 -524
rect 388 -560 444 -524
rect 480 -560 536 -524
rect 572 -560 590 -524
rect 0 -600 590 -560
<< nsubdiff >>
rect 0 3330 554 3360
rect 0 3294 18 3330
rect 54 3294 110 3330
rect 146 3294 202 3330
rect 238 3294 294 3330
rect 330 3294 386 3330
rect 422 3294 478 3330
rect 514 3294 554 3330
rect 0 3238 554 3294
rect 0 3202 18 3238
rect 54 3202 110 3238
rect 146 3202 202 3238
rect 238 3202 294 3238
rect 330 3202 386 3238
rect 422 3202 478 3238
rect 514 3202 554 3238
rect 0 3160 554 3202
<< psubdiffcont >>
rect 76 -468 112 -432
rect 168 -468 204 -432
rect 260 -468 296 -432
rect 352 -468 388 -432
rect 444 -468 480 -432
rect 536 -468 572 -432
rect 76 -560 112 -524
rect 168 -560 204 -524
rect 260 -560 296 -524
rect 352 -560 388 -524
rect 444 -560 480 -524
rect 536 -560 572 -524
<< nsubdiffcont >>
rect 18 3294 54 3330
rect 110 3294 146 3330
rect 202 3294 238 3330
rect 294 3294 330 3330
rect 386 3294 422 3330
rect 478 3294 514 3330
rect 662 3294 698 3330
rect 18 3202 54 3238
rect 110 3202 146 3238
rect 202 3202 238 3238
rect 294 3202 330 3238
rect 386 3202 422 3238
rect 478 3202 514 3238
<< poly >>
rect 0 1076 66 1092
rect 0 1042 16 1076
rect 50 1056 66 1076
rect 218 1056 248 1166
rect 50 1044 492 1056
rect 50 1042 66 1044
rect 0 1026 66 1042
rect 188 1014 366 1044
<< polycont >>
rect 16 1042 50 1076
<< locali >>
rect -36 3330 590 3346
rect -36 3294 18 3330
rect 54 3294 110 3330
rect 146 3294 202 3330
rect 238 3294 294 3330
rect 330 3294 386 3330
rect 422 3294 478 3330
rect 514 3294 590 3330
rect -36 3238 590 3294
rect -36 3202 18 3238
rect 54 3202 110 3238
rect 146 3202 202 3238
rect 238 3202 294 3238
rect 330 3202 386 3238
rect 422 3202 478 3238
rect 514 3202 590 3238
rect -36 3174 590 3202
rect 172 1596 206 3174
rect 0 1076 66 1092
rect 0 1042 16 1076
rect 50 1042 66 1076
rect 260 1066 294 1188
rect 488 1076 554 1092
rect 488 1066 504 1076
rect 0 1026 66 1042
rect 108 1042 504 1066
rect 538 1042 554 1076
rect 108 1026 554 1042
rect 108 992 142 1026
rect 412 992 446 1026
rect 12 -416 46 84
rect 204 -416 238 84
rect 316 -416 350 84
rect 508 -416 542 84
rect 0 -432 590 -416
rect 0 -468 76 -432
rect 112 -468 168 -432
rect 204 -468 260 -432
rect 296 -468 352 -432
rect 388 -468 444 -432
rect 480 -468 536 -432
rect 572 -468 590 -432
rect 0 -524 590 -468
rect 0 -560 76 -524
rect 112 -560 168 -524
rect 204 -560 260 -524
rect 296 -560 352 -524
rect 388 -560 444 -524
rect 480 -560 536 -524
rect 572 -560 590 -524
rect 0 -584 590 -560
<< viali >>
rect 18 3294 54 3330
rect 110 3294 146 3330
rect 202 3294 238 3330
rect 294 3294 330 3330
rect 386 3294 422 3330
rect 478 3294 514 3330
rect 18 3202 54 3238
rect 110 3202 146 3238
rect 202 3202 238 3238
rect 294 3202 330 3238
rect 386 3202 422 3238
rect 478 3202 514 3238
rect 16 1042 50 1076
rect 504 1042 538 1076
rect 76 -468 112 -432
rect 168 -468 204 -432
rect 260 -468 296 -432
rect 352 -468 388 -432
rect 444 -468 480 -432
rect 536 -468 572 -432
rect 76 -560 112 -524
rect 168 -560 204 -524
rect 260 -560 296 -524
rect 352 -560 388 -524
rect 444 -560 480 -524
rect 536 -560 572 -524
<< metal1 >>
rect -36 3330 590 3346
rect -36 3294 18 3330
rect 54 3294 110 3330
rect 146 3294 202 3330
rect 238 3294 294 3330
rect 330 3294 386 3330
rect 422 3294 478 3330
rect 514 3294 590 3330
rect -36 3238 590 3294
rect -36 3202 18 3238
rect 54 3202 110 3238
rect 146 3202 202 3238
rect 238 3202 294 3238
rect 330 3202 386 3238
rect 422 3202 478 3238
rect 514 3202 590 3238
rect -36 3174 590 3202
rect 0 1076 66 1092
rect 0 1042 16 1076
rect 50 1042 66 1076
rect 0 1026 66 1042
rect 488 1076 554 1092
rect 488 1042 504 1076
rect 538 1042 554 1076
rect 488 1026 554 1042
rect 0 -432 590 -416
rect 0 -468 76 -432
rect 112 -468 168 -432
rect 204 -468 260 -432
rect 296 -468 352 -432
rect 388 -468 444 -432
rect 480 -468 536 -432
rect 572 -468 590 -432
rect 0 -524 590 -468
rect 0 -560 76 -524
rect 112 -560 168 -524
rect 204 -560 260 -524
rect 296 -560 352 -524
rect 388 -560 444 -524
rect 480 -560 536 -524
rect 572 -560 590 -524
rect 0 -584 590 -560
use sky130_fd_pr__nfet_01v8_QQ9VTX  sky130_fd_pr__nfet_01v8_QQ9VTX_0
timestamp 1755919380
transform 1 0 125 0 1 538
box -125 -476 125 506
use sky130_fd_pr__nfet_01v8_QQ9VTX  sky130_fd_pr__nfet_01v8_QQ9VTX_1
timestamp 1755919380
transform 1 0 429 0 1 538
box -125 -476 125 506
use sky130_fd_pr__pfet_01v8_UCB5V5  sky130_fd_pr__pfet_01v8_UCB5V5_0
timestamp 1755919380
transform 1 0 233 0 1 1392
box -109 -262 109 262
<< end >>
