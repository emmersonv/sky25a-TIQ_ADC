magic
tech sky130A
timestamp 1755723063
<< nwell >>
rect 100 428 118 446
rect 139 428 157 446
rect 231 428 249 446
rect 270 428 288 446
rect 100 382 118 400
rect 139 382 157 400
rect 231 382 249 400
rect 270 382 288 400
rect 100 -64 118 -46
rect 139 -64 157 -46
rect 231 -64 249 -46
rect 270 -64 288 -46
rect 100 -110 118 -92
rect 139 -110 157 -92
rect 231 -110 249 -92
rect 270 -110 288 -92
rect 100 -557 118 -539
rect 139 -557 157 -539
rect 231 -557 249 -539
rect 270 -557 288 -539
rect 100 -603 118 -585
rect 139 -603 157 -585
rect 231 -603 249 -585
rect 270 -603 288 -585
rect 100 -1049 118 -1031
rect 139 -1049 157 -1031
rect 231 -1049 249 -1031
rect 270 -1049 288 -1031
rect 100 -1095 118 -1077
rect 139 -1095 157 -1077
rect 231 -1095 249 -1077
rect 270 -1095 288 -1077
rect 100 -1541 118 -1523
rect 139 -1541 157 -1523
rect 231 -1541 249 -1523
rect 270 -1541 288 -1523
rect 100 -1587 118 -1569
rect 139 -1587 157 -1569
rect 231 -1587 249 -1569
rect 270 -1587 288 -1569
rect 100 -2033 118 -2015
rect 139 -2033 157 -2015
rect 231 -2033 249 -2015
rect 270 -2033 288 -2015
rect 100 -2079 118 -2061
rect 139 -2079 157 -2061
rect 231 -2079 249 -2061
rect 270 -2079 288 -2061
rect 100 -2525 118 -2507
rect 139 -2525 157 -2507
rect 231 -2525 249 -2507
rect 270 -2525 288 -2507
rect 100 -2571 118 -2553
rect 139 -2571 157 -2553
rect 231 -2571 249 -2553
rect 270 -2571 288 -2553
<< psubdiff >>
rect 0 8 393 92
rect 0 -484 393 -400
rect -1 -977 394 -892
rect 0 -1470 393 -1385
rect 0 -1961 393 -1877
rect 0 -2453 393 -2368
rect 0 -2945 393 -2861
<< nsubdiffcont >>
rect 100 428 118 446
rect 139 428 157 446
rect 231 428 249 446
rect 270 428 288 446
rect 100 382 118 400
rect 139 382 157 400
rect 231 382 249 400
rect 270 382 288 400
rect 100 -64 118 -46
rect 139 -64 157 -46
rect 231 -64 249 -46
rect 270 -64 288 -46
rect 100 -110 118 -92
rect 139 -110 157 -92
rect 231 -110 249 -92
rect 270 -110 288 -92
rect 100 -557 118 -539
rect 139 -557 157 -539
rect 231 -557 249 -539
rect 270 -557 288 -539
rect 100 -603 118 -585
rect 139 -603 157 -585
rect 231 -603 249 -585
rect 270 -603 288 -585
rect 100 -1049 118 -1031
rect 139 -1049 157 -1031
rect 231 -1049 249 -1031
rect 270 -1049 288 -1031
rect 100 -1095 118 -1077
rect 139 -1095 157 -1077
rect 231 -1095 249 -1077
rect 270 -1095 288 -1077
rect 100 -1541 118 -1523
rect 139 -1541 157 -1523
rect 231 -1541 249 -1523
rect 270 -1541 288 -1523
rect 100 -1587 118 -1569
rect 139 -1587 157 -1569
rect 231 -1587 249 -1569
rect 270 -1587 288 -1569
rect 100 -2033 118 -2015
rect 139 -2033 157 -2015
rect 231 -2033 249 -2015
rect 270 -2033 288 -2015
rect 100 -2079 118 -2061
rect 139 -2079 157 -2061
rect 231 -2079 249 -2061
rect 270 -2079 288 -2061
rect 100 -2525 118 -2507
rect 139 -2525 157 -2507
rect 231 -2525 249 -2507
rect 270 -2525 288 -2507
rect 100 -2571 118 -2553
rect 139 -2571 157 -2553
rect 231 -2571 249 -2553
rect 270 -2571 288 -2553
<< locali >>
rect 0 182 33 216
rect 369 188 393 208
rect 0 8 393 92
rect 0 -310 33 -276
rect 369 -304 393 -284
rect 0 -484 393 -400
rect 0 -803 33 -769
rect 369 -797 393 -777
rect -1 -977 394 -892
rect 0 -1295 33 -1261
rect 369 -1289 393 -1269
rect 0 -1470 393 -1385
rect 0 -1787 33 -1753
rect 369 -1781 393 -1761
rect 0 -1961 393 -1877
rect 0 -2279 33 -2245
rect 369 -2273 393 -2253
rect 0 -2453 393 -2368
rect 0 -2771 33 -2737
rect 369 -2765 393 -2745
rect 0 -2945 393 -2861
<< viali >>
rect 100 428 118 446
rect 139 428 157 446
rect 231 428 249 446
rect 270 428 288 446
rect 100 382 118 400
rect 139 382 157 400
rect 231 382 249 400
rect 270 382 288 400
rect 100 -64 118 -46
rect 139 -64 157 -46
rect 231 -64 249 -46
rect 270 -64 288 -46
rect 100 -110 118 -92
rect 139 -110 157 -92
rect 231 -110 249 -92
rect 270 -110 288 -92
rect 100 -557 118 -539
rect 139 -557 157 -539
rect 231 -557 249 -539
rect 270 -557 288 -539
rect 100 -603 118 -585
rect 139 -603 157 -585
rect 231 -603 249 -585
rect 270 -603 288 -585
rect 100 -1049 118 -1031
rect 139 -1049 157 -1031
rect 231 -1049 249 -1031
rect 270 -1049 288 -1031
rect 100 -1095 118 -1077
rect 139 -1095 157 -1077
rect 231 -1095 249 -1077
rect 270 -1095 288 -1077
rect 100 -1541 118 -1523
rect 139 -1541 157 -1523
rect 231 -1541 249 -1523
rect 270 -1541 288 -1523
rect 100 -1587 118 -1569
rect 139 -1587 157 -1569
rect 231 -1587 249 -1569
rect 270 -1587 288 -1569
rect 100 -2033 118 -2015
rect 139 -2033 157 -2015
rect 231 -2033 249 -2015
rect 270 -2033 288 -2015
rect 100 -2079 118 -2061
rect 139 -2079 157 -2061
rect 231 -2079 249 -2061
rect 270 -2079 288 -2061
rect 100 -2525 118 -2507
rect 139 -2525 157 -2507
rect 231 -2525 249 -2507
rect 270 -2525 288 -2507
rect 100 -2571 118 -2553
rect 139 -2571 157 -2553
rect 231 -2571 249 -2553
rect 270 -2571 288 -2553
<< metal1 >>
rect 0 446 394 454
rect 0 428 100 446
rect 118 428 139 446
rect 157 428 231 446
rect 249 428 270 446
rect 288 428 394 446
rect 0 400 394 428
rect 0 382 100 400
rect 118 382 139 400
rect 157 382 231 400
rect 249 382 270 400
rect 288 382 394 400
rect 0 368 394 382
rect 0 8 393 92
rect 1 -46 395 -37
rect 1 -64 100 -46
rect 118 -64 139 -46
rect 157 -64 231 -46
rect 249 -64 270 -46
rect 288 -64 395 -46
rect 1 -92 395 -64
rect 1 -110 100 -92
rect 118 -110 139 -92
rect 157 -110 231 -92
rect 249 -110 270 -92
rect 288 -110 395 -92
rect 1 -123 395 -110
rect 0 -484 393 -400
rect 0 -539 394 -531
rect 0 -557 100 -539
rect 118 -557 139 -539
rect 157 -557 231 -539
rect 249 -557 270 -539
rect 288 -557 394 -539
rect 0 -585 394 -557
rect 0 -603 100 -585
rect 118 -603 139 -585
rect 157 -603 231 -585
rect 249 -603 270 -585
rect 288 -603 394 -585
rect 0 -617 394 -603
rect -1 -977 394 -892
rect 0 -1031 394 -1023
rect 0 -1049 100 -1031
rect 118 -1049 139 -1031
rect 157 -1049 231 -1031
rect 249 -1049 270 -1031
rect 288 -1049 394 -1031
rect 0 -1077 394 -1049
rect 0 -1095 100 -1077
rect 118 -1095 139 -1077
rect 157 -1095 231 -1077
rect 249 -1095 270 -1077
rect 288 -1095 394 -1077
rect 0 -1109 394 -1095
rect 0 -1470 393 -1385
rect 0 -1523 394 -1515
rect 0 -1541 100 -1523
rect 118 -1541 139 -1523
rect 157 -1541 231 -1523
rect 249 -1541 270 -1523
rect 288 -1541 394 -1523
rect 0 -1569 394 -1541
rect 0 -1587 100 -1569
rect 118 -1587 139 -1569
rect 157 -1587 231 -1569
rect 249 -1587 270 -1569
rect 288 -1587 394 -1569
rect 0 -1601 394 -1587
rect 0 -1961 393 -1877
rect 0 -2015 394 -2007
rect 0 -2033 100 -2015
rect 118 -2033 139 -2015
rect 157 -2033 231 -2015
rect 249 -2033 270 -2015
rect 288 -2033 394 -2015
rect 0 -2061 394 -2033
rect 0 -2079 100 -2061
rect 118 -2079 139 -2061
rect 157 -2079 231 -2061
rect 249 -2079 270 -2061
rect 288 -2079 394 -2061
rect 0 -2093 394 -2079
rect 0 -2453 393 -2368
rect 0 -2507 394 -2499
rect 0 -2525 100 -2507
rect 118 -2525 139 -2507
rect 157 -2525 231 -2507
rect 249 -2525 270 -2507
rect 288 -2525 394 -2507
rect 0 -2553 394 -2525
rect 0 -2571 100 -2553
rect 118 -2571 139 -2553
rect 157 -2571 231 -2553
rect 249 -2571 270 -2553
rect 288 -2571 394 -2553
rect 0 -2585 394 -2571
rect 0 -2945 393 -2861
use gain_stage  gain_stage_0
timestamp 1754266322
transform 1 0 0 0 1 0
box 0 0 393 479
use gain_stage  gain_stage_1
timestamp 1754266322
transform 1 0 0 0 1 -492
box 0 0 393 479
use gain_stage  gain_stage_2
timestamp 1754266322
transform 1 0 0 0 1 -985
box 0 0 393 479
use gain_stage  gain_stage_3
timestamp 1754266322
transform 1 0 0 0 1 -1477
box 0 0 393 479
use gain_stage  gain_stage_4
timestamp 1754266322
transform 1 0 0 0 1 -1969
box 0 0 393 479
use gain_stage  gain_stage_5
timestamp 1754266322
transform 1 0 0 0 1 -2461
box 0 0 393 479
use gain_stage  gain_stage_6
timestamp 1754266322
transform 1 0 0 0 1 -2953
box 0 0 393 479
<< end >>
