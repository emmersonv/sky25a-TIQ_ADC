magic
tech sky130A
magscale 1 2
timestamp 1755919380
<< error_s >>
rect -592 216 -576 366
rect -540 216 -322 470
rect -592 198 -322 216
rect -540 188 -436 198
<< nwell >>
rect -540 2312 678 2540
rect -512 2286 648 2312
rect -492 2254 -458 2286
rect -300 2254 -266 2286
rect 4 2254 38 2286
rect 196 2254 230 2286
rect 404 2254 438 2286
rect 596 2254 630 2286
rect -592 198 -576 216
<< psubdiff >>
rect -638 -1288 730 -1256
rect -638 -1324 -608 -1288
rect -572 -1324 -516 -1288
rect -480 -1324 -424 -1288
rect -388 -1324 -332 -1288
rect -296 -1324 -240 -1288
rect -204 -1324 -148 -1288
rect -112 -1324 -56 -1288
rect -20 -1324 36 -1288
rect 72 -1324 128 -1288
rect 164 -1324 220 -1288
rect 256 -1324 312 -1288
rect 348 -1324 404 -1288
rect 440 -1324 496 -1288
rect 532 -1324 588 -1288
rect 624 -1324 680 -1288
rect 716 -1324 730 -1288
rect -638 -1380 730 -1324
rect -638 -1416 -608 -1380
rect -572 -1416 -516 -1380
rect -480 -1416 -424 -1380
rect -388 -1416 -332 -1380
rect -296 -1416 -240 -1380
rect -204 -1416 -148 -1380
rect -112 -1416 -56 -1380
rect -20 -1416 36 -1380
rect 72 -1416 128 -1380
rect 164 -1416 220 -1380
rect 256 -1416 312 -1380
rect 348 -1416 404 -1380
rect 440 -1416 496 -1380
rect 532 -1416 588 -1380
rect 624 -1416 680 -1380
rect 716 -1416 730 -1380
rect -638 -1456 730 -1416
<< nsubdiff >>
rect -504 2474 642 2504
rect -504 2438 -482 2474
rect -446 2438 -390 2474
rect -354 2438 -298 2474
rect -262 2438 -206 2474
rect -170 2438 -114 2474
rect -78 2438 -22 2474
rect 14 2438 70 2474
rect 106 2438 162 2474
rect 198 2438 254 2474
rect 290 2438 346 2474
rect 382 2438 438 2474
rect 474 2438 530 2474
rect 566 2438 642 2474
rect -504 2382 642 2438
rect -504 2346 -482 2382
rect -446 2346 -390 2382
rect -354 2346 -298 2382
rect -262 2346 -206 2382
rect -170 2346 -114 2382
rect -78 2346 -22 2382
rect 14 2346 70 2382
rect 106 2346 162 2382
rect 198 2346 254 2382
rect 290 2346 346 2382
rect 382 2346 438 2382
rect 474 2346 530 2382
rect 566 2346 642 2382
rect -504 2304 642 2346
<< psubdiffcont >>
rect -608 -1324 -572 -1288
rect -516 -1324 -480 -1288
rect -424 -1324 -388 -1288
rect -332 -1324 -296 -1288
rect -240 -1324 -204 -1288
rect -148 -1324 -112 -1288
rect -56 -1324 -20 -1288
rect 36 -1324 72 -1288
rect 128 -1324 164 -1288
rect 220 -1324 256 -1288
rect 312 -1324 348 -1288
rect 404 -1324 440 -1288
rect 496 -1324 532 -1288
rect 588 -1324 624 -1288
rect 680 -1324 716 -1288
rect -608 -1416 -572 -1380
rect -516 -1416 -480 -1380
rect -424 -1416 -388 -1380
rect -332 -1416 -296 -1380
rect -240 -1416 -204 -1380
rect -148 -1416 -112 -1380
rect -56 -1416 -20 -1380
rect 36 -1416 72 -1380
rect 128 -1416 164 -1380
rect 220 -1416 256 -1380
rect 312 -1416 348 -1380
rect 404 -1416 440 -1380
rect 496 -1416 532 -1380
rect 588 -1416 624 -1380
rect 680 -1416 716 -1380
<< nsubdiffcont >>
rect -482 2438 -446 2474
rect -390 2438 -354 2474
rect -298 2438 -262 2474
rect -206 2438 -170 2474
rect -114 2438 -78 2474
rect -22 2438 14 2474
rect 70 2438 106 2474
rect 162 2438 198 2474
rect 254 2438 290 2474
rect 346 2438 382 2474
rect 438 2438 474 2474
rect 530 2438 566 2474
rect -482 2346 -446 2382
rect -390 2346 -354 2382
rect -298 2346 -262 2382
rect -206 2346 -170 2382
rect -114 2346 -78 2382
rect -22 2346 14 2382
rect 70 2346 106 2382
rect 162 2346 198 2382
rect 254 2346 290 2382
rect 346 2346 382 2382
rect 438 2346 474 2382
rect 530 2346 566 2382
<< poly >>
rect -592 220 -526 236
rect -592 186 -576 220
rect -542 200 -526 220
rect -542 194 -394 200
rect -220 194 -42 224
rect 180 194 358 224
rect -542 186 580 194
rect -592 170 580 186
rect 58 146 88 170
<< polycont >>
rect -576 186 -542 220
<< locali >>
rect -592 2474 730 2490
rect -592 2438 -574 2474
rect -538 2438 -482 2474
rect -446 2438 -390 2474
rect -354 2438 -298 2474
rect -262 2438 -206 2474
rect -170 2438 -114 2474
rect -78 2438 -22 2474
rect 14 2438 70 2474
rect 106 2438 162 2474
rect 198 2438 254 2474
rect 290 2438 346 2474
rect 382 2438 438 2474
rect 474 2438 530 2474
rect 566 2438 622 2474
rect 658 2438 730 2474
rect -592 2382 730 2438
rect -592 2346 -574 2382
rect -538 2346 -482 2382
rect -446 2346 -390 2382
rect -354 2346 -298 2382
rect -262 2346 -206 2382
rect -170 2346 -114 2382
rect -78 2346 -22 2382
rect 14 2346 70 2382
rect 106 2346 162 2382
rect 198 2346 254 2382
rect 290 2346 346 2382
rect 382 2346 438 2382
rect 474 2346 530 2382
rect 566 2346 622 2382
rect 658 2346 730 2382
rect -592 2318 730 2346
rect -492 2254 -458 2318
rect -300 2254 -266 2318
rect 4 2254 38 2318
rect 196 2254 230 2318
rect 404 2254 438 2318
rect 596 2254 630 2318
rect -592 220 -526 236
rect -592 186 -576 220
rect -542 186 -526 220
rect -592 170 -526 186
rect -396 208 -362 246
rect -204 208 -170 246
rect -92 212 -58 246
rect 100 212 134 246
rect 308 212 342 246
rect 500 212 534 246
rect 664 222 730 238
rect 664 212 680 222
rect -92 208 680 212
rect -396 188 680 208
rect 714 188 730 222
rect -396 172 730 188
rect -396 170 -54 172
rect 100 124 134 172
rect 12 -1272 46 22
rect -638 -1288 730 -1272
rect -638 -1324 -608 -1288
rect -572 -1324 -516 -1288
rect -480 -1324 -424 -1288
rect -388 -1324 -332 -1288
rect -296 -1324 -240 -1288
rect -204 -1324 -148 -1288
rect -112 -1324 -56 -1288
rect -20 -1324 36 -1288
rect 72 -1324 128 -1288
rect 164 -1324 220 -1288
rect 256 -1324 312 -1288
rect 348 -1324 404 -1288
rect 440 -1324 496 -1288
rect 532 -1324 588 -1288
rect 624 -1324 680 -1288
rect 716 -1324 730 -1288
rect -638 -1380 730 -1324
rect -638 -1416 -608 -1380
rect -572 -1416 -516 -1380
rect -480 -1416 -424 -1380
rect -388 -1416 -332 -1380
rect -296 -1416 -240 -1380
rect -204 -1416 -148 -1380
rect -112 -1416 -56 -1380
rect -20 -1416 36 -1380
rect 72 -1416 128 -1380
rect 164 -1416 220 -1380
rect 256 -1416 312 -1380
rect 348 -1416 404 -1380
rect 440 -1416 496 -1380
rect 532 -1416 588 -1380
rect 624 -1416 680 -1380
rect 716 -1416 730 -1380
rect -638 -1440 730 -1416
<< viali >>
rect -574 2438 -538 2474
rect -482 2438 -446 2474
rect -390 2438 -354 2474
rect -298 2438 -262 2474
rect -206 2438 -170 2474
rect -114 2438 -78 2474
rect -22 2438 14 2474
rect 70 2438 106 2474
rect 162 2438 198 2474
rect 254 2438 290 2474
rect 346 2438 382 2474
rect 438 2438 474 2474
rect 530 2438 566 2474
rect 622 2438 658 2474
rect -574 2346 -538 2382
rect -482 2346 -446 2382
rect -390 2346 -354 2382
rect -298 2346 -262 2382
rect -206 2346 -170 2382
rect -114 2346 -78 2382
rect -22 2346 14 2382
rect 70 2346 106 2382
rect 162 2346 198 2382
rect 254 2346 290 2382
rect 346 2346 382 2382
rect 438 2346 474 2382
rect 530 2346 566 2382
rect 622 2346 658 2382
rect -576 186 -542 220
rect 680 188 714 222
rect -608 -1324 -572 -1288
rect -516 -1324 -480 -1288
rect -424 -1324 -388 -1288
rect -332 -1324 -296 -1288
rect -240 -1324 -204 -1288
rect -148 -1324 -112 -1288
rect -56 -1324 -20 -1288
rect 36 -1324 72 -1288
rect 128 -1324 164 -1288
rect 220 -1324 256 -1288
rect 312 -1324 348 -1288
rect 404 -1324 440 -1288
rect 496 -1324 532 -1288
rect 588 -1324 624 -1288
rect 680 -1324 716 -1288
rect -608 -1416 -572 -1380
rect -516 -1416 -480 -1380
rect -424 -1416 -388 -1380
rect -332 -1416 -296 -1380
rect -240 -1416 -204 -1380
rect -148 -1416 -112 -1380
rect -56 -1416 -20 -1380
rect 36 -1416 72 -1380
rect 128 -1416 164 -1380
rect 220 -1416 256 -1380
rect 312 -1416 348 -1380
rect 404 -1416 440 -1380
rect 496 -1416 532 -1380
rect 588 -1416 624 -1380
rect 680 -1416 716 -1380
<< metal1 >>
rect -592 2474 730 2490
rect -592 2438 -574 2474
rect -538 2438 -482 2474
rect -446 2438 -390 2474
rect -354 2438 -298 2474
rect -262 2438 -206 2474
rect -170 2438 -114 2474
rect -78 2438 -22 2474
rect 14 2438 70 2474
rect 106 2438 162 2474
rect 198 2438 254 2474
rect 290 2438 346 2474
rect 382 2438 438 2474
rect 474 2438 530 2474
rect 566 2438 622 2474
rect 658 2438 730 2474
rect -592 2382 730 2438
rect -592 2346 -574 2382
rect -538 2346 -482 2382
rect -446 2346 -390 2382
rect -354 2346 -298 2382
rect -262 2346 -206 2382
rect -170 2346 -114 2382
rect -78 2346 -22 2382
rect 14 2346 70 2382
rect 106 2346 162 2382
rect 198 2346 254 2382
rect 290 2346 346 2382
rect 382 2346 438 2382
rect 474 2346 530 2382
rect 566 2346 622 2382
rect 658 2346 730 2382
rect -592 2318 730 2346
rect -592 220 -526 236
rect -592 186 -576 220
rect -542 186 -526 220
rect -592 170 -526 186
rect 664 222 730 238
rect 664 188 680 222
rect 714 188 730 222
rect 664 172 730 188
rect -638 -1288 730 -1272
rect -638 -1324 -608 -1288
rect -572 -1324 -516 -1288
rect -480 -1324 -424 -1288
rect -388 -1324 -332 -1288
rect -296 -1324 -240 -1288
rect -204 -1324 -148 -1288
rect -112 -1324 -56 -1288
rect -20 -1324 36 -1288
rect 72 -1324 128 -1288
rect 164 -1324 220 -1288
rect 256 -1324 312 -1288
rect 348 -1324 404 -1288
rect 440 -1324 496 -1288
rect 532 -1324 588 -1288
rect 624 -1324 680 -1288
rect 716 -1324 730 -1288
rect -638 -1380 730 -1324
rect -638 -1416 -608 -1380
rect -572 -1416 -516 -1380
rect -480 -1416 -424 -1380
rect -388 -1416 -332 -1380
rect -296 -1416 -240 -1380
rect -204 -1416 -148 -1380
rect -112 -1416 -56 -1380
rect -20 -1416 36 -1380
rect 72 -1416 128 -1380
rect 164 -1416 220 -1380
rect 256 -1416 312 -1380
rect 348 -1416 404 -1380
rect 440 -1416 496 -1380
rect 532 -1416 588 -1380
rect 624 -1416 680 -1380
rect 716 -1416 730 -1380
rect -638 -1440 730 -1416
use sky130_fd_pr__nfet_01v8_PD6K7A  sky130_fd_pr__nfet_01v8_PD6K7A_0
timestamp 1755919380
transform 1 0 73 0 1 73
box -73 -73 73 73
use sky130_fd_pr__pfet_01v8_WGHLR5  sky130_fd_pr__pfet_01v8_WGHLR5_0
timestamp 1755919380
transform 1 0 -331 0 1 1250
box -209 -1062 209 1062
use sky130_fd_pr__pfet_01v8_WGHLR5  sky130_fd_pr__pfet_01v8_WGHLR5_1
timestamp 1755919380
transform 1 0 69 0 1 1250
box -209 -1062 209 1062
use sky130_fd_pr__pfet_01v8_WGHLR5  sky130_fd_pr__pfet_01v8_WGHLR5_2
timestamp 1755919380
transform 1 0 469 0 1 1250
box -209 -1062 209 1062
<< end >>
