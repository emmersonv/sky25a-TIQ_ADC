magic
tech sky130A
timestamp 1755911681
<< polycont >>
rect 370 3143 387 3161
rect 370 2651 387 2669
rect 370 2158 387 2176
rect 370 1666 387 1684
rect 370 1174 387 1192
rect 370 682 387 700
rect 370 190 387 208
<< locali >>
rect 362 3161 395 3169
rect 2 3141 26 3161
rect 362 3143 370 3161
rect 387 3143 395 3161
rect 362 3135 395 3143
rect 448 2908 532 2941
rect 448 2890 460 2908
rect 478 2890 532 2908
rect 362 2669 395 2677
rect 2 2649 26 2669
rect 362 2651 370 2669
rect 387 2651 395 2669
rect 362 2643 395 2651
rect 362 2176 395 2184
rect 2 2156 26 2176
rect 362 2158 370 2176
rect 387 2158 395 2176
rect 362 2150 395 2158
rect 362 1684 395 1692
rect 2 1664 26 1684
rect 362 1666 370 1684
rect 387 1666 395 1684
rect 362 1658 395 1666
rect 362 1192 395 1200
rect 2 1172 26 1192
rect 362 1174 370 1192
rect 387 1174 395 1192
rect 362 1166 395 1174
rect 362 700 395 708
rect 2 680 26 700
rect 362 682 370 700
rect 387 682 395 700
rect 362 674 395 682
rect 448 379 532 2890
rect 2327 894 2413 2941
rect 2327 876 2387 894
rect 2405 876 2413 894
rect 2327 380 2413 876
rect 362 208 395 216
rect 2 188 26 208
rect 362 190 370 208
rect 387 190 395 208
rect 362 182 395 190
<< viali >>
rect 370 3143 387 3161
rect 460 2890 478 2908
rect 370 2651 387 2669
rect 370 2158 387 2176
rect 370 1666 387 1684
rect 370 1174 387 1192
rect 370 682 387 700
rect 2387 876 2405 894
rect 370 190 387 208
<< metal1 >>
rect -130 3321 2 3407
rect 395 3321 2413 3409
rect -130 2916 -55 3321
rect 362 3166 395 3169
rect 362 3139 365 3166
rect 392 3139 395 3166
rect 362 3135 395 3139
rect 395 2962 541 3046
rect 440 2941 541 2962
rect -130 2830 2 2916
rect 448 2908 532 2941
rect 448 2890 460 2908
rect 478 2890 532 2908
rect -130 2422 -55 2830
rect 362 2674 395 2677
rect 362 2647 365 2674
rect 392 2647 395 2674
rect 362 2643 395 2647
rect 448 2553 532 2890
rect 395 2469 532 2553
rect -130 2336 2 2422
rect -130 1930 -55 2336
rect 362 2180 395 2184
rect 362 2153 365 2180
rect 392 2153 395 2180
rect 362 2150 395 2153
rect 448 2061 532 2469
rect 396 1977 532 2061
rect -130 1844 3 1930
rect -130 1438 -55 1844
rect 362 1689 395 1692
rect 362 1662 365 1689
rect 392 1662 395 1689
rect 362 1658 395 1662
rect 448 1568 532 1977
rect 395 1484 532 1568
rect -130 1352 2 1438
rect -130 946 -55 1352
rect 362 1197 395 1200
rect 362 1170 365 1197
rect 392 1170 395 1197
rect 362 1166 395 1170
rect 448 1077 532 1484
rect 395 993 532 1077
rect -130 860 2 946
rect -130 454 -55 860
rect 362 705 395 708
rect 362 678 365 705
rect 392 678 395 705
rect 362 674 395 678
rect 448 585 532 993
rect 395 501 532 585
rect -130 368 1 454
rect 362 213 395 216
rect 362 186 365 213
rect 392 186 395 213
rect 362 182 395 186
rect 448 92 532 501
rect 2327 894 2413 3321
rect 2327 876 2387 894
rect 2405 876 2413 894
rect 2327 380 2413 876
rect 395 8 532 92
<< via1 >>
rect 365 3161 392 3166
rect 365 3143 370 3161
rect 370 3143 387 3161
rect 387 3143 392 3161
rect 365 3139 392 3143
rect 365 2669 392 2674
rect 365 2651 370 2669
rect 370 2651 387 2669
rect 387 2651 392 2669
rect 365 2647 392 2651
rect 365 2176 392 2180
rect 365 2158 370 2176
rect 370 2158 387 2176
rect 387 2158 392 2176
rect 365 2153 392 2158
rect 365 1684 392 1689
rect 365 1666 370 1684
rect 370 1666 387 1684
rect 387 1666 392 1684
rect 365 1662 392 1666
rect 365 1192 392 1197
rect 365 1174 370 1192
rect 370 1174 387 1192
rect 387 1174 392 1192
rect 365 1170 392 1174
rect 365 700 392 705
rect 365 682 370 700
rect 370 682 387 700
rect 387 682 392 700
rect 365 678 392 682
rect 365 208 392 213
rect 365 190 370 208
rect 370 190 387 208
rect 387 190 392 208
rect 365 186 392 190
<< metal2 >>
rect 362 3166 1232 3169
rect 362 3139 365 3166
rect 392 3139 1232 3166
rect 362 3135 1232 3139
rect 362 2674 1185 2677
rect 362 2647 365 2674
rect 392 2647 1185 2674
rect 362 2643 1185 2647
rect 1152 2223 1185 2643
rect 1199 2527 1232 3135
rect 1199 2494 1286 2527
rect 1152 2190 1286 2223
rect 362 2180 1138 2184
rect 362 2153 365 2180
rect 392 2153 1138 2180
rect 362 2150 1138 2153
rect 1105 1919 1138 2150
rect 1105 1886 1286 1919
rect 362 1689 1286 1695
rect 362 1662 365 1689
rect 392 1662 1286 1689
rect 362 1658 395 1662
rect 1199 1440 1253 1473
rect 1199 1200 1232 1440
rect 362 1197 1232 1200
rect 362 1170 365 1197
rect 392 1170 1232 1197
rect 362 1166 1232 1170
rect 1199 1058 1253 1091
rect 1199 708 1232 1058
rect 1301 1016 1318 2915
rect 362 705 1232 708
rect 362 678 365 705
rect 392 678 1232 705
rect 362 674 1232 678
rect 1254 216 1287 380
rect 362 213 1287 216
rect 362 186 365 213
rect 392 186 1287 213
rect 362 182 1287 186
use gain_stage_7  gain_stage_7_0
timestamp 1755723063
transform -1 0 395 0 1 2953
box -1 -2953 395 479
use tiq_adc_7  tiq_adc_7_0
timestamp 1755723063
transform 1 0 440 0 1 380
box 0 0 1998 2561
<< labels >>
rlabel metal1 1184 3321 1266 3409 1 VDPWR
port 1 n
rlabel metal1 448 8 529 86 5 VGND
port 2 s
rlabel metal2 1301 1779 1318 1802 3 Vin
port 3 e
rlabel locali 5 3145 18 3157 7 t0
port 4 w
rlabel locali 6 2653 19 2665 7 t1
port 5 w
rlabel locali 5 2159 18 2171 7 t2
port 6 w
rlabel locali 5 1668 18 1680 7 t3
port 7 w
rlabel locali 5 1176 18 1188 7 t4
port 8 w
rlabel locali 5 684 18 696 7 t5
port 9 w
rlabel locali 4 192 17 204 7 t6
port 10 w
<< end >>
