magic
tech sky130A
magscale 1 2
timestamp 1756008383
<< error_s >>
rect -142 2996 290 3128
rect -142 2960 -36 2996
rect 26 2960 122 2996
rect 0 2760 280 2960
rect 552 2760 554 2960
rect 588 2724 590 2996
<< nwell >>
rect -36 2960 588 2996
rect -36 2760 26 2960
rect 122 2760 588 2960
rect -36 2172 588 2760
rect -36 656 590 2172
<< pwell >>
rect -26 -1026 580 -774
<< psubdiff >>
rect 0 -833 554 -800
rect 0 -867 21 -833
rect 55 -867 113 -833
rect 147 -867 205 -833
rect 239 -867 297 -833
rect 331 -867 389 -833
rect 423 -867 481 -833
rect 515 -867 554 -833
rect 0 -925 554 -867
rect 0 -959 21 -925
rect 55 -959 113 -925
rect 147 -959 205 -925
rect 239 -959 297 -925
rect 331 -959 389 -925
rect 423 -959 481 -925
rect 515 -959 554 -925
rect 0 -1000 554 -959
<< nsubdiff >>
rect 0 2760 26 2960
rect 122 2929 554 2960
rect 122 2895 147 2929
rect 181 2895 239 2929
rect 273 2895 331 2929
rect 365 2895 423 2929
rect 457 2895 554 2929
rect 122 2837 554 2895
rect 122 2803 147 2837
rect 181 2803 239 2837
rect 273 2803 331 2837
rect 365 2803 423 2837
rect 457 2803 554 2837
rect 122 2760 554 2803
<< psubdiffcont >>
rect 21 -867 55 -833
rect 113 -867 147 -833
rect 205 -867 239 -833
rect 297 -867 331 -833
rect 389 -867 423 -833
rect 481 -867 515 -833
rect 21 -959 55 -925
rect 113 -959 147 -925
rect 205 -959 239 -925
rect 297 -959 331 -925
rect 389 -959 423 -925
rect 481 -959 515 -925
<< nsubdiffcont >>
rect 147 2895 181 2929
rect 239 2895 273 2929
rect 331 2895 365 2929
rect 423 2895 457 2929
rect 147 2803 181 2837
rect 239 2803 273 2837
rect 331 2803 365 2837
rect 423 2803 457 2837
<< poly >>
rect 0 676 66 692
rect 0 642 16 676
rect 50 656 66 676
rect 218 656 248 692
rect 50 644 492 656
rect 50 642 66 644
rect 0 626 66 642
rect 188 614 366 644
<< polycont >>
rect 16 642 50 676
<< locali >>
rect -36 2774 26 2946
rect 122 2929 590 2946
rect 122 2895 147 2929
rect 181 2895 239 2929
rect 273 2895 331 2929
rect 365 2895 423 2929
rect 457 2895 515 2929
rect 549 2895 590 2929
rect 122 2837 590 2895
rect 122 2803 147 2837
rect 181 2803 239 2837
rect 273 2803 331 2837
rect 365 2803 423 2837
rect 457 2803 515 2837
rect 549 2803 590 2837
rect 122 2774 590 2803
rect 172 2106 206 2774
rect 0 676 66 692
rect 0 642 16 676
rect 50 642 66 676
rect 260 666 294 714
rect 488 676 554 692
rect 488 666 504 676
rect 0 626 66 642
rect 108 642 504 666
rect 538 642 554 676
rect 108 626 554 642
rect 108 576 142 626
rect 412 592 446 626
rect 12 -816 46 84
rect 204 -816 238 84
rect 316 -816 350 84
rect 508 -816 542 84
rect -36 -833 588 -816
rect -36 -867 21 -833
rect 55 -867 113 -833
rect 147 -867 205 -833
rect 239 -867 297 -833
rect 331 -867 389 -833
rect 423 -867 481 -833
rect 515 -867 588 -833
rect -36 -925 588 -867
rect -36 -959 21 -925
rect 55 -959 113 -925
rect 147 -959 205 -925
rect 239 -959 297 -925
rect 331 -959 389 -925
rect 423 -959 481 -925
rect 515 -959 588 -925
rect -36 -984 588 -959
<< viali >>
rect 147 2895 181 2929
rect 239 2895 273 2929
rect 331 2895 365 2929
rect 423 2895 457 2929
rect 515 2895 549 2929
rect 147 2803 181 2837
rect 239 2803 273 2837
rect 331 2803 365 2837
rect 423 2803 457 2837
rect 515 2803 549 2837
rect 16 642 50 676
rect 504 642 538 676
rect 21 -867 55 -833
rect 113 -867 147 -833
rect 205 -867 239 -833
rect 297 -867 331 -833
rect 389 -867 423 -833
rect 481 -867 515 -833
rect 21 -959 55 -925
rect 113 -959 147 -925
rect 205 -959 239 -925
rect 297 -959 331 -925
rect 389 -959 423 -925
rect 481 -959 515 -925
<< metal1 >>
rect -36 2774 26 2946
rect 122 2929 590 2946
rect 122 2895 147 2929
rect 181 2895 239 2929
rect 273 2895 331 2929
rect 365 2895 423 2929
rect 457 2895 515 2929
rect 549 2895 590 2929
rect 122 2837 590 2895
rect 122 2803 147 2837
rect 181 2803 239 2837
rect 273 2803 331 2837
rect 365 2803 423 2837
rect 457 2803 515 2837
rect 549 2803 590 2837
rect 122 2774 590 2803
rect 0 676 66 692
rect 0 642 16 676
rect 50 642 66 676
rect 0 626 66 642
rect 488 676 554 692
rect 488 642 504 676
rect 538 642 554 676
rect 488 626 554 642
rect -36 -833 588 -816
rect -36 -867 21 -833
rect 55 -867 113 -833
rect 147 -867 205 -833
rect 239 -867 297 -833
rect 331 -867 389 -833
rect 423 -867 481 -833
rect 515 -867 588 -833
rect -36 -925 588 -867
rect -36 -959 21 -925
rect 55 -959 113 -925
rect 147 -959 205 -925
rect 239 -959 297 -925
rect 331 -959 389 -925
rect 423 -959 481 -925
rect 515 -959 588 -925
rect -36 -984 588 -959
use sky130_fd_pr__nfet_01v8_V2VUT3  sky130_fd_pr__nfet_01v8_V2VUT3_0
timestamp 1756008383
transform 1 0 125 0 1 338
box -151 -276 151 306
use sky130_fd_pr__nfet_01v8_V2VUT3  sky130_fd_pr__nfet_01v8_V2VUT3_1
timestamp 1756008383
transform 1 0 429 0 1 338
box -151 -276 151 306
use sky130_fd_pr__pfet_01v8_VGLYR5  sky130_fd_pr__pfet_01v8_VGLYR5_0
timestamp 1756008383
transform 1 0 233 0 1 1418
box -109 -762 109 762
<< end >>
