magic
tech sky130A
magscale 1 2
timestamp 1756008383
<< nwell >>
rect -161 -812 161 812
<< pmos >>
rect -63 -750 -33 750
rect 33 -750 63 750
<< pdiff >>
rect -125 731 -63 750
rect -125 697 -113 731
rect -79 697 -63 731
rect -125 663 -63 697
rect -125 629 -113 663
rect -79 629 -63 663
rect -125 595 -63 629
rect -125 561 -113 595
rect -79 561 -63 595
rect -125 527 -63 561
rect -125 493 -113 527
rect -79 493 -63 527
rect -125 459 -63 493
rect -125 425 -113 459
rect -79 425 -63 459
rect -125 391 -63 425
rect -125 357 -113 391
rect -79 357 -63 391
rect -125 323 -63 357
rect -125 289 -113 323
rect -79 289 -63 323
rect -125 255 -63 289
rect -125 221 -113 255
rect -79 221 -63 255
rect -125 187 -63 221
rect -125 153 -113 187
rect -79 153 -63 187
rect -125 119 -63 153
rect -125 85 -113 119
rect -79 85 -63 119
rect -125 51 -63 85
rect -125 17 -113 51
rect -79 17 -63 51
rect -125 -17 -63 17
rect -125 -51 -113 -17
rect -79 -51 -63 -17
rect -125 -85 -63 -51
rect -125 -119 -113 -85
rect -79 -119 -63 -85
rect -125 -153 -63 -119
rect -125 -187 -113 -153
rect -79 -187 -63 -153
rect -125 -221 -63 -187
rect -125 -255 -113 -221
rect -79 -255 -63 -221
rect -125 -289 -63 -255
rect -125 -323 -113 -289
rect -79 -323 -63 -289
rect -125 -357 -63 -323
rect -125 -391 -113 -357
rect -79 -391 -63 -357
rect -125 -425 -63 -391
rect -125 -459 -113 -425
rect -79 -459 -63 -425
rect -125 -493 -63 -459
rect -125 -527 -113 -493
rect -79 -527 -63 -493
rect -125 -561 -63 -527
rect -125 -595 -113 -561
rect -79 -595 -63 -561
rect -125 -629 -63 -595
rect -125 -663 -113 -629
rect -79 -663 -63 -629
rect -125 -697 -63 -663
rect -125 -731 -113 -697
rect -79 -731 -63 -697
rect -125 -750 -63 -731
rect -33 731 33 750
rect -33 697 -17 731
rect 17 697 33 731
rect -33 663 33 697
rect -33 629 -17 663
rect 17 629 33 663
rect -33 595 33 629
rect -33 561 -17 595
rect 17 561 33 595
rect -33 527 33 561
rect -33 493 -17 527
rect 17 493 33 527
rect -33 459 33 493
rect -33 425 -17 459
rect 17 425 33 459
rect -33 391 33 425
rect -33 357 -17 391
rect 17 357 33 391
rect -33 323 33 357
rect -33 289 -17 323
rect 17 289 33 323
rect -33 255 33 289
rect -33 221 -17 255
rect 17 221 33 255
rect -33 187 33 221
rect -33 153 -17 187
rect 17 153 33 187
rect -33 119 33 153
rect -33 85 -17 119
rect 17 85 33 119
rect -33 51 33 85
rect -33 17 -17 51
rect 17 17 33 51
rect -33 -17 33 17
rect -33 -51 -17 -17
rect 17 -51 33 -17
rect -33 -85 33 -51
rect -33 -119 -17 -85
rect 17 -119 33 -85
rect -33 -153 33 -119
rect -33 -187 -17 -153
rect 17 -187 33 -153
rect -33 -221 33 -187
rect -33 -255 -17 -221
rect 17 -255 33 -221
rect -33 -289 33 -255
rect -33 -323 -17 -289
rect 17 -323 33 -289
rect -33 -357 33 -323
rect -33 -391 -17 -357
rect 17 -391 33 -357
rect -33 -425 33 -391
rect -33 -459 -17 -425
rect 17 -459 33 -425
rect -33 -493 33 -459
rect -33 -527 -17 -493
rect 17 -527 33 -493
rect -33 -561 33 -527
rect -33 -595 -17 -561
rect 17 -595 33 -561
rect -33 -629 33 -595
rect -33 -663 -17 -629
rect 17 -663 33 -629
rect -33 -697 33 -663
rect -33 -731 -17 -697
rect 17 -731 33 -697
rect -33 -750 33 -731
rect 63 731 125 750
rect 63 697 79 731
rect 113 697 125 731
rect 63 663 125 697
rect 63 629 79 663
rect 113 629 125 663
rect 63 595 125 629
rect 63 561 79 595
rect 113 561 125 595
rect 63 527 125 561
rect 63 493 79 527
rect 113 493 125 527
rect 63 459 125 493
rect 63 425 79 459
rect 113 425 125 459
rect 63 391 125 425
rect 63 357 79 391
rect 113 357 125 391
rect 63 323 125 357
rect 63 289 79 323
rect 113 289 125 323
rect 63 255 125 289
rect 63 221 79 255
rect 113 221 125 255
rect 63 187 125 221
rect 63 153 79 187
rect 113 153 125 187
rect 63 119 125 153
rect 63 85 79 119
rect 113 85 125 119
rect 63 51 125 85
rect 63 17 79 51
rect 113 17 125 51
rect 63 -17 125 17
rect 63 -51 79 -17
rect 113 -51 125 -17
rect 63 -85 125 -51
rect 63 -119 79 -85
rect 113 -119 125 -85
rect 63 -153 125 -119
rect 63 -187 79 -153
rect 113 -187 125 -153
rect 63 -221 125 -187
rect 63 -255 79 -221
rect 113 -255 125 -221
rect 63 -289 125 -255
rect 63 -323 79 -289
rect 113 -323 125 -289
rect 63 -357 125 -323
rect 63 -391 79 -357
rect 113 -391 125 -357
rect 63 -425 125 -391
rect 63 -459 79 -425
rect 113 -459 125 -425
rect 63 -493 125 -459
rect 63 -527 79 -493
rect 113 -527 125 -493
rect 63 -561 125 -527
rect 63 -595 79 -561
rect 113 -595 125 -561
rect 63 -629 125 -595
rect 63 -663 79 -629
rect 113 -663 125 -629
rect 63 -697 125 -663
rect 63 -731 79 -697
rect 113 -731 125 -697
rect 63 -750 125 -731
<< pdiffc >>
rect -113 697 -79 731
rect -113 629 -79 663
rect -113 561 -79 595
rect -113 493 -79 527
rect -113 425 -79 459
rect -113 357 -79 391
rect -113 289 -79 323
rect -113 221 -79 255
rect -113 153 -79 187
rect -113 85 -79 119
rect -113 17 -79 51
rect -113 -51 -79 -17
rect -113 -119 -79 -85
rect -113 -187 -79 -153
rect -113 -255 -79 -221
rect -113 -323 -79 -289
rect -113 -391 -79 -357
rect -113 -459 -79 -425
rect -113 -527 -79 -493
rect -113 -595 -79 -561
rect -113 -663 -79 -629
rect -113 -731 -79 -697
rect -17 697 17 731
rect -17 629 17 663
rect -17 561 17 595
rect -17 493 17 527
rect -17 425 17 459
rect -17 357 17 391
rect -17 289 17 323
rect -17 221 17 255
rect -17 153 17 187
rect -17 85 17 119
rect -17 17 17 51
rect -17 -51 17 -17
rect -17 -119 17 -85
rect -17 -187 17 -153
rect -17 -255 17 -221
rect -17 -323 17 -289
rect -17 -391 17 -357
rect -17 -459 17 -425
rect -17 -527 17 -493
rect -17 -595 17 -561
rect -17 -663 17 -629
rect -17 -731 17 -697
rect 79 697 113 731
rect 79 629 113 663
rect 79 561 113 595
rect 79 493 113 527
rect 79 425 113 459
rect 79 357 113 391
rect 79 289 113 323
rect 79 221 113 255
rect 79 153 113 187
rect 79 85 113 119
rect 79 17 113 51
rect 79 -51 113 -17
rect 79 -119 113 -85
rect 79 -187 113 -153
rect 79 -255 113 -221
rect 79 -323 113 -289
rect 79 -391 113 -357
rect 79 -459 113 -425
rect 79 -527 113 -493
rect 79 -595 113 -561
rect 79 -663 113 -629
rect 79 -731 113 -697
<< poly >>
rect -63 750 -33 780
rect 33 750 63 780
rect -63 -776 -33 -750
rect 33 -776 63 -750
rect -63 -806 63 -776
<< locali >>
rect -113 737 -79 754
rect -113 665 -79 697
rect -113 595 -79 629
rect -113 527 -79 559
rect -113 459 -79 487
rect -113 391 -79 415
rect -113 323 -79 343
rect -113 255 -79 271
rect -113 187 -79 199
rect -113 119 -79 127
rect -113 51 -79 55
rect -113 -55 -79 -51
rect -113 -127 -79 -119
rect -113 -199 -79 -187
rect -113 -271 -79 -255
rect -113 -343 -79 -323
rect -113 -415 -79 -391
rect -113 -487 -79 -459
rect -113 -559 -79 -527
rect -113 -629 -79 -595
rect -113 -697 -79 -665
rect -113 -754 -79 -737
rect -17 737 17 754
rect -17 665 17 697
rect -17 595 17 629
rect -17 527 17 559
rect -17 459 17 487
rect -17 391 17 415
rect -17 323 17 343
rect -17 255 17 271
rect -17 187 17 199
rect -17 119 17 127
rect -17 51 17 55
rect -17 -55 17 -51
rect -17 -127 17 -119
rect -17 -199 17 -187
rect -17 -271 17 -255
rect -17 -343 17 -323
rect -17 -415 17 -391
rect -17 -487 17 -459
rect -17 -559 17 -527
rect -17 -629 17 -595
rect -17 -697 17 -665
rect -17 -754 17 -737
rect 79 737 113 754
rect 79 665 113 697
rect 79 595 113 629
rect 79 527 113 559
rect 79 459 113 487
rect 79 391 113 415
rect 79 323 113 343
rect 79 255 113 271
rect 79 187 113 199
rect 79 119 113 127
rect 79 51 113 55
rect 79 -55 113 -51
rect 79 -127 113 -119
rect 79 -199 113 -187
rect 79 -271 113 -255
rect 79 -343 113 -323
rect 79 -415 113 -391
rect 79 -487 113 -459
rect 79 -559 113 -527
rect 79 -629 113 -595
rect 79 -697 113 -665
rect 79 -754 113 -737
<< viali >>
rect -113 731 -79 737
rect -113 703 -79 731
rect -113 663 -79 665
rect -113 631 -79 663
rect -113 561 -79 593
rect -113 559 -79 561
rect -113 493 -79 521
rect -113 487 -79 493
rect -113 425 -79 449
rect -113 415 -79 425
rect -113 357 -79 377
rect -113 343 -79 357
rect -113 289 -79 305
rect -113 271 -79 289
rect -113 221 -79 233
rect -113 199 -79 221
rect -113 153 -79 161
rect -113 127 -79 153
rect -113 85 -79 89
rect -113 55 -79 85
rect -113 -17 -79 17
rect -113 -85 -79 -55
rect -113 -89 -79 -85
rect -113 -153 -79 -127
rect -113 -161 -79 -153
rect -113 -221 -79 -199
rect -113 -233 -79 -221
rect -113 -289 -79 -271
rect -113 -305 -79 -289
rect -113 -357 -79 -343
rect -113 -377 -79 -357
rect -113 -425 -79 -415
rect -113 -449 -79 -425
rect -113 -493 -79 -487
rect -113 -521 -79 -493
rect -113 -561 -79 -559
rect -113 -593 -79 -561
rect -113 -663 -79 -631
rect -113 -665 -79 -663
rect -113 -731 -79 -703
rect -113 -737 -79 -731
rect -17 731 17 737
rect -17 703 17 731
rect -17 663 17 665
rect -17 631 17 663
rect -17 561 17 593
rect -17 559 17 561
rect -17 493 17 521
rect -17 487 17 493
rect -17 425 17 449
rect -17 415 17 425
rect -17 357 17 377
rect -17 343 17 357
rect -17 289 17 305
rect -17 271 17 289
rect -17 221 17 233
rect -17 199 17 221
rect -17 153 17 161
rect -17 127 17 153
rect -17 85 17 89
rect -17 55 17 85
rect -17 -17 17 17
rect -17 -85 17 -55
rect -17 -89 17 -85
rect -17 -153 17 -127
rect -17 -161 17 -153
rect -17 -221 17 -199
rect -17 -233 17 -221
rect -17 -289 17 -271
rect -17 -305 17 -289
rect -17 -357 17 -343
rect -17 -377 17 -357
rect -17 -425 17 -415
rect -17 -449 17 -425
rect -17 -493 17 -487
rect -17 -521 17 -493
rect -17 -561 17 -559
rect -17 -593 17 -561
rect -17 -663 17 -631
rect -17 -665 17 -663
rect -17 -731 17 -703
rect -17 -737 17 -731
rect 79 731 113 737
rect 79 703 113 731
rect 79 663 113 665
rect 79 631 113 663
rect 79 561 113 593
rect 79 559 113 561
rect 79 493 113 521
rect 79 487 113 493
rect 79 425 113 449
rect 79 415 113 425
rect 79 357 113 377
rect 79 343 113 357
rect 79 289 113 305
rect 79 271 113 289
rect 79 221 113 233
rect 79 199 113 221
rect 79 153 113 161
rect 79 127 113 153
rect 79 85 113 89
rect 79 55 113 85
rect 79 -17 113 17
rect 79 -85 113 -55
rect 79 -89 113 -85
rect 79 -153 113 -127
rect 79 -161 113 -153
rect 79 -221 113 -199
rect 79 -233 113 -221
rect 79 -289 113 -271
rect 79 -305 113 -289
rect 79 -357 113 -343
rect 79 -377 113 -357
rect 79 -425 113 -415
rect 79 -449 113 -425
rect 79 -493 113 -487
rect 79 -521 113 -493
rect 79 -561 113 -559
rect 79 -593 113 -561
rect 79 -663 113 -631
rect 79 -665 113 -663
rect 79 -731 113 -703
rect 79 -737 113 -731
<< metal1 >>
rect -119 737 -73 750
rect -119 703 -113 737
rect -79 703 -73 737
rect -119 665 -73 703
rect -119 631 -113 665
rect -79 631 -73 665
rect -119 593 -73 631
rect -119 559 -113 593
rect -79 559 -73 593
rect -119 521 -73 559
rect -119 487 -113 521
rect -79 487 -73 521
rect -119 449 -73 487
rect -119 415 -113 449
rect -79 415 -73 449
rect -119 377 -73 415
rect -119 343 -113 377
rect -79 343 -73 377
rect -119 305 -73 343
rect -119 271 -113 305
rect -79 271 -73 305
rect -119 233 -73 271
rect -119 199 -113 233
rect -79 199 -73 233
rect -119 161 -73 199
rect -119 127 -113 161
rect -79 127 -73 161
rect -119 89 -73 127
rect -119 55 -113 89
rect -79 55 -73 89
rect -119 17 -73 55
rect -119 -17 -113 17
rect -79 -17 -73 17
rect -119 -55 -73 -17
rect -119 -89 -113 -55
rect -79 -89 -73 -55
rect -119 -127 -73 -89
rect -119 -161 -113 -127
rect -79 -161 -73 -127
rect -119 -199 -73 -161
rect -119 -233 -113 -199
rect -79 -233 -73 -199
rect -119 -271 -73 -233
rect -119 -305 -113 -271
rect -79 -305 -73 -271
rect -119 -343 -73 -305
rect -119 -377 -113 -343
rect -79 -377 -73 -343
rect -119 -415 -73 -377
rect -119 -449 -113 -415
rect -79 -449 -73 -415
rect -119 -487 -73 -449
rect -119 -521 -113 -487
rect -79 -521 -73 -487
rect -119 -559 -73 -521
rect -119 -593 -113 -559
rect -79 -593 -73 -559
rect -119 -631 -73 -593
rect -119 -665 -113 -631
rect -79 -665 -73 -631
rect -119 -703 -73 -665
rect -119 -737 -113 -703
rect -79 -737 -73 -703
rect -119 -750 -73 -737
rect -23 737 23 750
rect -23 703 -17 737
rect 17 703 23 737
rect -23 665 23 703
rect -23 631 -17 665
rect 17 631 23 665
rect -23 593 23 631
rect -23 559 -17 593
rect 17 559 23 593
rect -23 521 23 559
rect -23 487 -17 521
rect 17 487 23 521
rect -23 449 23 487
rect -23 415 -17 449
rect 17 415 23 449
rect -23 377 23 415
rect -23 343 -17 377
rect 17 343 23 377
rect -23 305 23 343
rect -23 271 -17 305
rect 17 271 23 305
rect -23 233 23 271
rect -23 199 -17 233
rect 17 199 23 233
rect -23 161 23 199
rect -23 127 -17 161
rect 17 127 23 161
rect -23 89 23 127
rect -23 55 -17 89
rect 17 55 23 89
rect -23 17 23 55
rect -23 -17 -17 17
rect 17 -17 23 17
rect -23 -55 23 -17
rect -23 -89 -17 -55
rect 17 -89 23 -55
rect -23 -127 23 -89
rect -23 -161 -17 -127
rect 17 -161 23 -127
rect -23 -199 23 -161
rect -23 -233 -17 -199
rect 17 -233 23 -199
rect -23 -271 23 -233
rect -23 -305 -17 -271
rect 17 -305 23 -271
rect -23 -343 23 -305
rect -23 -377 -17 -343
rect 17 -377 23 -343
rect -23 -415 23 -377
rect -23 -449 -17 -415
rect 17 -449 23 -415
rect -23 -487 23 -449
rect -23 -521 -17 -487
rect 17 -521 23 -487
rect -23 -559 23 -521
rect -23 -593 -17 -559
rect 17 -593 23 -559
rect -23 -631 23 -593
rect -23 -665 -17 -631
rect 17 -665 23 -631
rect -23 -703 23 -665
rect -23 -737 -17 -703
rect 17 -737 23 -703
rect -23 -750 23 -737
rect 73 737 119 750
rect 73 703 79 737
rect 113 703 119 737
rect 73 665 119 703
rect 73 631 79 665
rect 113 631 119 665
rect 73 593 119 631
rect 73 559 79 593
rect 113 559 119 593
rect 73 521 119 559
rect 73 487 79 521
rect 113 487 119 521
rect 73 449 119 487
rect 73 415 79 449
rect 113 415 119 449
rect 73 377 119 415
rect 73 343 79 377
rect 113 343 119 377
rect 73 305 119 343
rect 73 271 79 305
rect 113 271 119 305
rect 73 233 119 271
rect 73 199 79 233
rect 113 199 119 233
rect 73 161 119 199
rect 73 127 79 161
rect 113 127 119 161
rect 73 89 119 127
rect 73 55 79 89
rect 113 55 119 89
rect 73 17 119 55
rect 73 -17 79 17
rect 113 -17 119 17
rect 73 -55 119 -17
rect 73 -89 79 -55
rect 113 -89 119 -55
rect 73 -127 119 -89
rect 73 -161 79 -127
rect 113 -161 119 -127
rect 73 -199 119 -161
rect 73 -233 79 -199
rect 113 -233 119 -199
rect 73 -271 119 -233
rect 73 -305 79 -271
rect 113 -305 119 -271
rect 73 -343 119 -305
rect 73 -377 79 -343
rect 113 -377 119 -343
rect 73 -415 119 -377
rect 73 -449 79 -415
rect 113 -449 119 -415
rect 73 -487 119 -449
rect 73 -521 79 -487
rect 113 -521 119 -487
rect 73 -559 119 -521
rect 73 -593 79 -559
rect 113 -593 119 -559
rect 73 -631 119 -593
rect 73 -665 79 -631
rect 113 -665 119 -631
rect 73 -703 119 -665
rect 73 -737 79 -703
rect 113 -737 119 -703
rect 73 -750 119 -737
<< end >>
