magic
tech sky130A
magscale 1 2
timestamp 1756008383
<< error_p >>
rect -36 3346 590 3396
rect 0 3324 554 3346
rect 0 3310 36 3324
rect 518 3310 554 3324
rect 0 3196 36 3210
rect 518 3196 554 3210
rect 0 3174 554 3196
rect -36 3160 590 3174
rect -36 3124 172 3160
rect 206 3124 590 3160
rect 206 2914 340 3124
<< error_s >>
rect 206 1654 340 2914
<< nwell >>
rect 0 3346 554 3360
rect -36 3174 590 3346
rect 0 3160 554 3174
rect 172 1646 206 3160
rect -36 1130 590 1646
<< pwell >>
rect -26 -626 616 -374
<< psubdiff >>
rect 0 -433 590 -400
rect 0 -467 77 -433
rect 111 -467 169 -433
rect 203 -467 261 -433
rect 295 -467 353 -433
rect 387 -467 445 -433
rect 479 -467 537 -433
rect 571 -467 590 -433
rect 0 -525 590 -467
rect 0 -559 77 -525
rect 111 -559 169 -525
rect 203 -559 261 -525
rect 295 -559 353 -525
rect 387 -559 445 -525
rect 479 -559 537 -525
rect 571 -559 590 -525
rect 0 -600 590 -559
<< nsubdiff >>
rect 0 3329 554 3360
rect 0 3295 19 3329
rect 53 3295 111 3329
rect 145 3295 203 3329
rect 237 3295 295 3329
rect 329 3295 387 3329
rect 421 3295 479 3329
rect 513 3295 554 3329
rect 0 3237 554 3295
rect 0 3203 19 3237
rect 53 3203 111 3237
rect 145 3203 203 3237
rect 237 3203 295 3237
rect 329 3203 387 3237
rect 421 3203 479 3237
rect 513 3203 554 3237
rect 0 3160 554 3203
<< psubdiffcont >>
rect 77 -467 111 -433
rect 169 -467 203 -433
rect 261 -467 295 -433
rect 353 -467 387 -433
rect 445 -467 479 -433
rect 537 -467 571 -433
rect 77 -559 111 -525
rect 169 -559 203 -525
rect 261 -559 295 -525
rect 353 -559 387 -525
rect 445 -559 479 -525
rect 537 -559 571 -525
<< nsubdiffcont >>
rect 19 3295 53 3329
rect 111 3295 145 3329
rect 203 3295 237 3329
rect 295 3295 329 3329
rect 387 3295 421 3329
rect 479 3295 513 3329
rect 19 3203 53 3237
rect 111 3203 145 3237
rect 203 3203 237 3237
rect 295 3203 329 3237
rect 387 3203 421 3237
rect 479 3203 513 3237
<< poly >>
rect 0 1076 66 1092
rect 0 1042 16 1076
rect 50 1056 66 1076
rect 218 1056 248 1166
rect 50 1044 492 1056
rect 50 1042 66 1044
rect 0 1026 66 1042
rect 188 1014 366 1044
<< polycont >>
rect 16 1042 50 1076
<< locali >>
rect -36 3329 590 3346
rect -36 3295 19 3329
rect 53 3295 111 3329
rect 145 3295 203 3329
rect 237 3295 295 3329
rect 329 3295 387 3329
rect 421 3295 479 3329
rect 513 3295 590 3329
rect -36 3237 590 3295
rect -36 3203 19 3237
rect 53 3203 111 3237
rect 145 3203 203 3237
rect 237 3203 295 3237
rect 329 3203 387 3237
rect 421 3203 479 3237
rect 513 3203 590 3237
rect -36 3174 590 3203
rect 172 1596 206 3174
rect 0 1076 66 1092
rect 0 1042 16 1076
rect 50 1042 66 1076
rect 260 1066 294 1188
rect 488 1076 554 1092
rect 488 1066 504 1076
rect 0 1026 66 1042
rect 108 1042 504 1066
rect 538 1042 554 1076
rect 108 1026 554 1042
rect 108 992 142 1026
rect 412 992 446 1026
rect 12 -416 46 84
rect 204 -416 238 84
rect 316 -416 350 84
rect 508 -416 542 84
rect 0 -433 590 -416
rect 0 -467 77 -433
rect 111 -467 169 -433
rect 203 -467 261 -433
rect 295 -467 353 -433
rect 387 -467 445 -433
rect 479 -467 537 -433
rect 571 -467 590 -433
rect 0 -525 590 -467
rect 0 -559 77 -525
rect 111 -559 169 -525
rect 203 -559 261 -525
rect 295 -559 353 -525
rect 387 -559 445 -525
rect 479 -559 537 -525
rect 571 -559 590 -525
rect 0 -584 590 -559
<< viali >>
rect 19 3295 53 3329
rect 111 3295 145 3329
rect 203 3295 237 3329
rect 295 3295 329 3329
rect 387 3295 421 3329
rect 479 3295 513 3329
rect 19 3203 53 3237
rect 111 3203 145 3237
rect 203 3203 237 3237
rect 295 3203 329 3237
rect 387 3203 421 3237
rect 479 3203 513 3237
rect 16 1042 50 1076
rect 504 1042 538 1076
rect 77 -467 111 -433
rect 169 -467 203 -433
rect 261 -467 295 -433
rect 353 -467 387 -433
rect 445 -467 479 -433
rect 537 -467 571 -433
rect 77 -559 111 -525
rect 169 -559 203 -525
rect 261 -559 295 -525
rect 353 -559 387 -525
rect 445 -559 479 -525
rect 537 -559 571 -525
<< metal1 >>
rect -36 3329 590 3346
rect -36 3295 19 3329
rect 53 3295 111 3329
rect 145 3295 203 3329
rect 237 3295 295 3329
rect 329 3295 387 3329
rect 421 3295 479 3329
rect 513 3295 590 3329
rect -36 3237 590 3295
rect -36 3203 19 3237
rect 53 3203 111 3237
rect 145 3203 203 3237
rect 237 3203 295 3237
rect 329 3203 387 3237
rect 421 3203 479 3237
rect 513 3203 590 3237
rect -36 3174 590 3203
rect 0 1076 66 1092
rect 0 1042 16 1076
rect 50 1042 66 1076
rect 0 1026 66 1042
rect 488 1076 554 1092
rect 488 1042 504 1076
rect 538 1042 554 1076
rect 488 1026 554 1042
rect 0 -433 590 -416
rect 0 -467 77 -433
rect 111 -467 169 -433
rect 203 -467 261 -433
rect 295 -467 353 -433
rect 387 -467 445 -433
rect 479 -467 537 -433
rect 571 -467 590 -433
rect 0 -525 590 -467
rect 0 -559 77 -525
rect 111 -559 169 -525
rect 203 -559 261 -525
rect 295 -559 353 -525
rect 387 -559 445 -525
rect 479 -559 537 -525
rect 571 -559 590 -525
rect 0 -584 590 -559
use sky130_fd_pr__nfet_01v8_QQ9VTX  sky130_fd_pr__nfet_01v8_QQ9VTX_0
timestamp 1756008383
transform 1 0 125 0 1 538
box -151 -476 151 506
use sky130_fd_pr__nfet_01v8_QQ9VTX  sky130_fd_pr__nfet_01v8_QQ9VTX_1
timestamp 1756008383
transform 1 0 429 0 1 538
box -151 -476 151 506
use sky130_fd_pr__pfet_01v8_UCB5V5  sky130_fd_pr__pfet_01v8_UCB5V5_0
timestamp 1756008383
transform 1 0 233 0 1 1392
box -109 -262 109 262
<< end >>
