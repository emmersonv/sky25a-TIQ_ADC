magic
tech sky130A
magscale 1 2
timestamp 1755911681
<< locali >>
rect 208 6320 274 6336
rect 208 6284 224 6320
rect 258 6284 274 6320
rect 208 6268 274 6284
rect 208 5334 274 5348
rect 208 5298 224 5334
rect 258 5298 274 5334
rect 208 5280 274 5298
rect 208 4350 274 4366
rect 208 4314 224 4350
rect 258 4314 274 4350
rect 208 4298 274 4314
rect 208 3366 274 3382
rect 208 3330 224 3366
rect 258 3330 274 3366
rect 208 3314 274 3330
rect 208 2382 274 2398
rect 208 2346 224 2382
rect 258 2346 274 2382
rect 208 2330 274 2346
rect 208 1396 274 1412
rect 208 1360 224 1396
rect 258 1360 274 1396
rect 208 1344 274 1360
rect 208 412 274 428
rect 208 376 224 412
rect 258 376 274 412
rect 208 360 274 376
<< viali >>
rect 224 6284 258 6320
rect 224 5298 258 5334
rect 224 4314 258 4350
rect 224 3330 258 3366
rect 224 2346 258 2382
rect 224 1360 258 1396
rect 224 376 258 412
<< metal1 >>
rect -130 6814 5082 6820
rect -3860 6806 5082 6814
rect -3860 6752 -3850 6806
rect -3796 6752 -3770 6806
rect -3716 6752 -3690 6806
rect -3636 6752 -3610 6806
rect -3556 6752 5082 6806
rect -3860 6726 5082 6752
rect -3860 6672 -3850 6726
rect -3796 6672 -3770 6726
rect -3716 6672 -3690 6726
rect -3636 6672 -3610 6726
rect -3556 6672 5082 6726
rect -3860 6640 5082 6672
rect -130 6638 5082 6640
rect 208 6330 274 6336
rect 208 6276 214 6330
rect 268 6276 274 6330
rect 208 6268 274 6276
rect 208 5342 274 5348
rect 208 5288 214 5342
rect 268 5288 274 5342
rect 208 5280 274 5288
rect 208 4360 274 4366
rect 208 4306 214 4360
rect 268 4306 274 4360
rect 208 4298 274 4306
rect 208 3376 274 3382
rect 208 3322 214 3376
rect 268 3322 274 3376
rect 208 3314 274 3322
rect 208 2392 274 2398
rect 208 2338 214 2392
rect 268 2338 274 2392
rect 208 2330 274 2338
rect 208 1406 274 1412
rect 208 1352 214 1406
rect 268 1352 274 1406
rect 208 1344 274 1352
rect 208 422 274 428
rect 208 368 214 422
rect 268 368 274 422
rect 208 360 274 368
rect -3200 156 1324 184
rect -3200 102 -3188 156
rect -3134 102 -3108 156
rect -3054 102 -3028 156
rect -2974 102 -2948 156
rect -2894 102 1324 156
rect -3200 76 1324 102
rect -3200 22 -3188 76
rect -3134 22 -3108 76
rect -3054 22 -3028 76
rect -2974 22 -2948 76
rect -2894 22 1324 76
rect -3200 16 1324 22
<< via1 >>
rect -3850 6752 -3796 6806
rect -3770 6752 -3716 6806
rect -3690 6752 -3636 6806
rect -3610 6752 -3556 6806
rect -3850 6672 -3796 6726
rect -3770 6672 -3716 6726
rect -3690 6672 -3636 6726
rect -3610 6672 -3556 6726
rect 214 6320 268 6330
rect 214 6284 224 6320
rect 224 6284 258 6320
rect 258 6284 268 6320
rect 214 6276 268 6284
rect 214 5334 268 5342
rect 214 5298 224 5334
rect 224 5298 258 5334
rect 258 5298 268 5334
rect 214 5288 268 5298
rect 214 4350 268 4360
rect 214 4314 224 4350
rect 224 4314 258 4350
rect 258 4314 268 4350
rect 214 4306 268 4314
rect 214 3366 268 3376
rect 214 3330 224 3366
rect 224 3330 258 3366
rect 258 3330 268 3366
rect 214 3322 268 3330
rect 214 2382 268 2392
rect 214 2346 224 2382
rect 224 2346 258 2382
rect 258 2346 268 2382
rect 214 2338 268 2346
rect 214 1396 268 1406
rect 214 1360 224 1396
rect 224 1360 258 1396
rect 258 1360 268 1396
rect 214 1352 268 1360
rect 214 412 268 422
rect 214 376 224 412
rect 224 376 258 412
rect 258 376 268 412
rect 214 368 268 376
rect -3188 102 -3134 156
rect -3108 102 -3054 156
rect -3028 102 -2974 156
rect -2948 102 -2894 156
rect -3188 22 -3134 76
rect -3108 22 -3054 76
rect -3028 22 -2974 76
rect -2948 22 -2894 76
<< metal2 >>
rect -260 6818 -192 6828
rect -3860 6808 -3540 6814
rect -3860 6752 -3850 6808
rect -3794 6752 -3770 6808
rect -3714 6752 -3690 6808
rect -3634 6752 -3610 6808
rect -3554 6752 -3540 6808
rect -3860 6728 -3540 6752
rect -3860 6672 -3850 6728
rect -3794 6672 -3770 6728
rect -3714 6672 -3690 6728
rect -3634 6672 -3610 6728
rect -3554 6672 -3540 6728
rect -3860 6640 -3540 6672
rect -260 6762 -254 6818
rect -198 6762 -192 6818
rect -260 6336 -192 6762
rect -260 6330 274 6336
rect -260 6276 214 6330
rect 268 6276 274 6330
rect -260 6268 274 6276
rect -238 5732 -170 5742
rect -238 5676 -232 5732
rect -176 5676 -170 5732
rect -238 5348 -170 5676
rect -238 5342 274 5348
rect -238 5288 214 5342
rect 268 5288 274 5342
rect -238 5280 274 5288
rect -238 4644 -170 4654
rect -238 4588 -232 4644
rect -176 4588 -170 4644
rect -238 4366 -170 4588
rect -238 4360 274 4366
rect -238 4306 214 4360
rect 268 4306 274 4360
rect -238 4298 274 4306
rect -238 3558 -170 3568
rect -238 3502 -232 3558
rect -176 3502 -170 3558
rect 2862 3506 2896 3664
rect -238 3382 -170 3502
rect -238 3376 274 3382
rect -238 3322 214 3376
rect 268 3322 274 3376
rect -238 3314 274 3322
rect -238 2462 -170 2472
rect -238 2406 -232 2462
rect -176 2406 -170 2462
rect -238 2398 -170 2406
rect -238 2392 274 2398
rect -238 2338 214 2392
rect 268 2338 274 2392
rect -238 2330 274 2338
rect -238 1406 274 1412
rect -238 1384 214 1406
rect -238 1328 -232 1384
rect -176 1352 214 1384
rect 268 1352 274 1406
rect -176 1344 274 1352
rect -176 1328 -170 1344
rect -238 1314 -170 1328
rect -3818 324 -3762 1016
rect -238 422 274 428
rect -238 368 214 422
rect 268 368 274 422
rect -238 360 274 368
rect -238 298 -170 360
rect -238 242 -232 298
rect -176 242 -170 298
rect -238 232 -170 242
rect -3200 158 -2880 184
rect -3200 102 -3188 158
rect -3132 102 -3108 158
rect -3052 102 -3028 158
rect -2972 102 -2948 158
rect -2892 102 -2880 158
rect -3200 78 -2880 102
rect -3200 22 -3188 78
rect -3132 22 -3108 78
rect -3052 22 -3028 78
rect -2972 22 -2948 78
rect -2892 22 -2880 78
rect -3200 16 -2880 22
<< via2 >>
rect -3850 6806 -3794 6808
rect -3850 6752 -3796 6806
rect -3796 6752 -3794 6806
rect -3770 6806 -3714 6808
rect -3770 6752 -3716 6806
rect -3716 6752 -3714 6806
rect -3690 6806 -3634 6808
rect -3690 6752 -3636 6806
rect -3636 6752 -3634 6806
rect -3610 6806 -3554 6808
rect -3610 6752 -3556 6806
rect -3556 6752 -3554 6806
rect -3850 6726 -3794 6728
rect -3850 6672 -3796 6726
rect -3796 6672 -3794 6726
rect -3770 6726 -3714 6728
rect -3770 6672 -3716 6726
rect -3716 6672 -3714 6726
rect -3690 6726 -3634 6728
rect -3690 6672 -3636 6726
rect -3636 6672 -3634 6726
rect -3610 6726 -3554 6728
rect -3610 6672 -3556 6726
rect -3556 6672 -3554 6726
rect -254 6762 -198 6818
rect -232 5676 -176 5732
rect -232 4588 -176 4644
rect -232 3502 -176 3558
rect -232 2406 -176 2462
rect -232 1328 -176 1384
rect -232 242 -176 298
rect -3188 156 -3132 158
rect -3188 102 -3134 156
rect -3134 102 -3132 156
rect -3108 156 -3052 158
rect -3108 102 -3054 156
rect -3054 102 -3052 156
rect -3028 156 -2972 158
rect -3028 102 -2974 156
rect -2974 102 -2972 156
rect -2948 156 -2892 158
rect -2948 102 -2894 156
rect -2894 102 -2892 156
rect -3188 76 -3132 78
rect -3188 22 -3134 76
rect -3134 22 -3132 76
rect -3108 76 -3052 78
rect -3108 22 -3054 76
rect -3054 22 -3052 76
rect -3028 76 -2972 78
rect -3028 22 -2974 76
rect -2974 22 -2972 76
rect -2948 76 -2892 78
rect -2948 22 -2894 76
rect -2894 22 -2892 76
<< metal3 >>
rect -276 6818 -178 6840
rect -3860 6812 -3540 6814
rect -3860 6748 -3854 6812
rect -3790 6748 -3774 6812
rect -3710 6748 -3694 6812
rect -3630 6748 -3614 6812
rect -3550 6748 -3540 6812
rect -3860 6732 -3540 6748
rect -276 6762 -254 6818
rect -198 6762 -178 6818
rect -276 6742 -178 6762
rect -3860 6668 -3854 6732
rect -3790 6668 -3774 6732
rect -3710 6668 -3694 6732
rect -3630 6668 -3614 6732
rect -3550 6668 -3540 6732
rect -3860 6640 -3540 6668
rect -7516 5916 -7116 6036
rect -254 5732 -156 5754
rect -254 5676 -232 5732
rect -176 5676 -156 5732
rect -254 5656 -156 5676
rect -254 4644 -156 4664
rect -254 4588 -232 4644
rect -176 4588 -156 4644
rect -254 4566 -156 4588
rect -7514 3468 -7114 3588
rect -254 3558 -156 3578
rect -254 3502 -232 3558
rect -176 3502 -156 3558
rect -254 3480 -156 3502
rect -256 2462 -158 2486
rect -256 2406 -232 2462
rect -176 2406 -158 2462
rect -256 2388 -158 2406
rect -254 1384 -156 1400
rect -254 1328 -232 1384
rect -176 1328 -156 1384
rect -254 1302 -156 1328
rect -7516 1020 -7116 1140
rect -256 298 -158 316
rect -256 242 -232 298
rect -176 242 -158 298
rect -256 218 -158 242
rect -3200 162 -2880 184
rect -3200 98 -3192 162
rect -3128 98 -3112 162
rect -3048 98 -3032 162
rect -2968 98 -2952 162
rect -2888 98 -2880 162
rect -3200 82 -2880 98
rect -3200 18 -3192 82
rect -3128 18 -3112 82
rect -3048 18 -3032 82
rect -2968 18 -2952 82
rect -2888 18 -2880 82
rect -3200 16 -2880 18
<< via3 >>
rect -3854 6808 -3790 6812
rect -3854 6752 -3850 6808
rect -3850 6752 -3794 6808
rect -3794 6752 -3790 6808
rect -3854 6748 -3790 6752
rect -3774 6808 -3710 6812
rect -3774 6752 -3770 6808
rect -3770 6752 -3714 6808
rect -3714 6752 -3710 6808
rect -3774 6748 -3710 6752
rect -3694 6808 -3630 6812
rect -3694 6752 -3690 6808
rect -3690 6752 -3634 6808
rect -3634 6752 -3630 6808
rect -3694 6748 -3630 6752
rect -3614 6808 -3550 6812
rect -3614 6752 -3610 6808
rect -3610 6752 -3554 6808
rect -3554 6752 -3550 6808
rect -3614 6748 -3550 6752
rect -3854 6728 -3790 6732
rect -3854 6672 -3850 6728
rect -3850 6672 -3794 6728
rect -3794 6672 -3790 6728
rect -3854 6668 -3790 6672
rect -3774 6728 -3710 6732
rect -3774 6672 -3770 6728
rect -3770 6672 -3714 6728
rect -3714 6672 -3710 6728
rect -3774 6668 -3710 6672
rect -3694 6728 -3630 6732
rect -3694 6672 -3690 6728
rect -3690 6672 -3634 6728
rect -3634 6672 -3630 6728
rect -3694 6668 -3630 6672
rect -3614 6728 -3550 6732
rect -3614 6672 -3610 6728
rect -3610 6672 -3554 6728
rect -3554 6672 -3550 6728
rect -3614 6668 -3550 6672
rect -3192 158 -3128 162
rect -3192 102 -3188 158
rect -3188 102 -3132 158
rect -3132 102 -3128 158
rect -3192 98 -3128 102
rect -3112 158 -3048 162
rect -3112 102 -3108 158
rect -3108 102 -3052 158
rect -3052 102 -3048 158
rect -3112 98 -3048 102
rect -3032 158 -2968 162
rect -3032 102 -3028 158
rect -3028 102 -2972 158
rect -2972 102 -2968 158
rect -3032 98 -2968 102
rect -2952 158 -2888 162
rect -2952 102 -2948 158
rect -2948 102 -2892 158
rect -2892 102 -2888 158
rect -2952 98 -2888 102
rect -3192 78 -3128 82
rect -3192 22 -3188 78
rect -3188 22 -3132 78
rect -3132 22 -3128 78
rect -3192 18 -3128 22
rect -3112 78 -3048 82
rect -3112 22 -3108 78
rect -3108 22 -3052 78
rect -3052 22 -3048 78
rect -3112 18 -3048 22
rect -3032 78 -2968 82
rect -3032 22 -3028 78
rect -3028 22 -2972 78
rect -2972 22 -2968 78
rect -3032 18 -2968 22
rect -2952 78 -2888 82
rect -2952 22 -2948 78
rect -2948 22 -2892 78
rect -2892 22 -2888 78
rect -2952 18 -2888 22
<< metal4 >>
rect -3860 6812 -3540 6814
rect -3860 6748 -3854 6812
rect -3790 6748 -3774 6812
rect -3710 6748 -3694 6812
rect -3630 6748 -3614 6812
rect -3550 6748 -3540 6812
rect -3860 6732 -3540 6748
rect -3860 6668 -3854 6732
rect -3790 6668 -3774 6732
rect -3710 6668 -3694 6732
rect -3630 6668 -3614 6732
rect -3550 6668 -3540 6732
rect -3860 6500 -3540 6668
rect -3200 162 -2880 420
rect -3200 98 -3192 162
rect -3128 98 -3112 162
rect -3048 98 -3032 162
rect -2968 98 -2952 162
rect -2888 98 -2880 162
rect -3200 82 -2880 98
rect -3200 18 -3192 82
rect -3128 18 -3112 82
rect -3048 18 -3032 82
rect -2968 18 -2952 82
rect -2888 18 -2880 82
rect -3200 16 -2880 18
use boosted_tiq_adc_7  boosted_tiq_adc_7_0
timestamp 1755911681
transform 1 0 260 0 1 0
box -260 0 4876 6864
use encoder  encoder_0
timestamp 1755737846
transform 1 0 -7516 0 1 -76
box 0 0 7471 6928
<< labels >>
rlabel metal1 -548 16 -380 184 5 VGND
port 1 s
rlabel metal1 -658 6640 -494 6814 1 VDPWR
port 2 n
rlabel metal2 2862 3506 2896 3664 3 Vin
port 3 e
rlabel metal3 -7516 1020 -7116 1140 7 o0
port 4 w
rlabel metal3 -7514 3468 -7114 3588 7 o1
port 5 w
rlabel metal3 -7516 5916 -7116 6036 7 o2
port 6 w
<< end >>
