magic
tech sky130A
magscale 1 2
timestamp 1756008383
<< pwell >>
rect -151 -476 151 476
<< nmos >>
rect -63 -450 -33 450
rect 33 -450 63 450
<< ndiff >>
rect -125 425 -63 450
rect -125 391 -113 425
rect -79 391 -63 425
rect -125 357 -63 391
rect -125 323 -113 357
rect -79 323 -63 357
rect -125 289 -63 323
rect -125 255 -113 289
rect -79 255 -63 289
rect -125 221 -63 255
rect -125 187 -113 221
rect -79 187 -63 221
rect -125 153 -63 187
rect -125 119 -113 153
rect -79 119 -63 153
rect -125 85 -63 119
rect -125 51 -113 85
rect -79 51 -63 85
rect -125 17 -63 51
rect -125 -17 -113 17
rect -79 -17 -63 17
rect -125 -51 -63 -17
rect -125 -85 -113 -51
rect -79 -85 -63 -51
rect -125 -119 -63 -85
rect -125 -153 -113 -119
rect -79 -153 -63 -119
rect -125 -187 -63 -153
rect -125 -221 -113 -187
rect -79 -221 -63 -187
rect -125 -255 -63 -221
rect -125 -289 -113 -255
rect -79 -289 -63 -255
rect -125 -323 -63 -289
rect -125 -357 -113 -323
rect -79 -357 -63 -323
rect -125 -391 -63 -357
rect -125 -425 -113 -391
rect -79 -425 -63 -391
rect -125 -450 -63 -425
rect -33 425 33 450
rect -33 391 -17 425
rect 17 391 33 425
rect -33 357 33 391
rect -33 323 -17 357
rect 17 323 33 357
rect -33 289 33 323
rect -33 255 -17 289
rect 17 255 33 289
rect -33 221 33 255
rect -33 187 -17 221
rect 17 187 33 221
rect -33 153 33 187
rect -33 119 -17 153
rect 17 119 33 153
rect -33 85 33 119
rect -33 51 -17 85
rect 17 51 33 85
rect -33 17 33 51
rect -33 -17 -17 17
rect 17 -17 33 17
rect -33 -51 33 -17
rect -33 -85 -17 -51
rect 17 -85 33 -51
rect -33 -119 33 -85
rect -33 -153 -17 -119
rect 17 -153 33 -119
rect -33 -187 33 -153
rect -33 -221 -17 -187
rect 17 -221 33 -187
rect -33 -255 33 -221
rect -33 -289 -17 -255
rect 17 -289 33 -255
rect -33 -323 33 -289
rect -33 -357 -17 -323
rect 17 -357 33 -323
rect -33 -391 33 -357
rect -33 -425 -17 -391
rect 17 -425 33 -391
rect -33 -450 33 -425
rect 63 425 125 450
rect 63 391 79 425
rect 113 391 125 425
rect 63 357 125 391
rect 63 323 79 357
rect 113 323 125 357
rect 63 289 125 323
rect 63 255 79 289
rect 113 255 125 289
rect 63 221 125 255
rect 63 187 79 221
rect 113 187 125 221
rect 63 153 125 187
rect 63 119 79 153
rect 113 119 125 153
rect 63 85 125 119
rect 63 51 79 85
rect 113 51 125 85
rect 63 17 125 51
rect 63 -17 79 17
rect 113 -17 125 17
rect 63 -51 125 -17
rect 63 -85 79 -51
rect 113 -85 125 -51
rect 63 -119 125 -85
rect 63 -153 79 -119
rect 113 -153 125 -119
rect 63 -187 125 -153
rect 63 -221 79 -187
rect 113 -221 125 -187
rect 63 -255 125 -221
rect 63 -289 79 -255
rect 113 -289 125 -255
rect 63 -323 125 -289
rect 63 -357 79 -323
rect 113 -357 125 -323
rect 63 -391 125 -357
rect 63 -425 79 -391
rect 113 -425 125 -391
rect 63 -450 125 -425
<< ndiffc >>
rect -113 391 -79 425
rect -113 323 -79 357
rect -113 255 -79 289
rect -113 187 -79 221
rect -113 119 -79 153
rect -113 51 -79 85
rect -113 -17 -79 17
rect -113 -85 -79 -51
rect -113 -153 -79 -119
rect -113 -221 -79 -187
rect -113 -289 -79 -255
rect -113 -357 -79 -323
rect -113 -425 -79 -391
rect -17 391 17 425
rect -17 323 17 357
rect -17 255 17 289
rect -17 187 17 221
rect -17 119 17 153
rect -17 51 17 85
rect -17 -17 17 17
rect -17 -85 17 -51
rect -17 -153 17 -119
rect -17 -221 17 -187
rect -17 -289 17 -255
rect -17 -357 17 -323
rect -17 -425 17 -391
rect 79 391 113 425
rect 79 323 113 357
rect 79 255 113 289
rect 79 187 113 221
rect 79 119 113 153
rect 79 51 113 85
rect 79 -17 113 17
rect 79 -85 113 -51
rect 79 -153 113 -119
rect 79 -221 113 -187
rect 79 -289 113 -255
rect 79 -357 113 -323
rect 79 -425 113 -391
<< poly >>
rect -63 476 63 506
rect -63 450 -33 476
rect 33 450 63 476
rect -63 -476 -33 -450
rect 33 -476 63 -450
<< locali >>
rect -113 425 -79 454
rect -113 357 -79 379
rect -113 289 -79 307
rect -113 221 -79 235
rect -113 153 -79 163
rect -113 85 -79 91
rect -113 17 -79 19
rect -113 -19 -79 -17
rect -113 -91 -79 -85
rect -113 -163 -79 -153
rect -113 -235 -79 -221
rect -113 -307 -79 -289
rect -113 -379 -79 -357
rect -113 -454 -79 -425
rect -17 425 17 454
rect -17 357 17 379
rect -17 289 17 307
rect -17 221 17 235
rect -17 153 17 163
rect -17 85 17 91
rect -17 17 17 19
rect -17 -19 17 -17
rect -17 -91 17 -85
rect -17 -163 17 -153
rect -17 -235 17 -221
rect -17 -307 17 -289
rect -17 -379 17 -357
rect -17 -454 17 -425
rect 79 425 113 454
rect 79 357 113 379
rect 79 289 113 307
rect 79 221 113 235
rect 79 153 113 163
rect 79 85 113 91
rect 79 17 113 19
rect 79 -19 113 -17
rect 79 -91 113 -85
rect 79 -163 113 -153
rect 79 -235 113 -221
rect 79 -307 113 -289
rect 79 -379 113 -357
rect 79 -454 113 -425
<< viali >>
rect -113 391 -79 413
rect -113 379 -79 391
rect -113 323 -79 341
rect -113 307 -79 323
rect -113 255 -79 269
rect -113 235 -79 255
rect -113 187 -79 197
rect -113 163 -79 187
rect -113 119 -79 125
rect -113 91 -79 119
rect -113 51 -79 53
rect -113 19 -79 51
rect -113 -51 -79 -19
rect -113 -53 -79 -51
rect -113 -119 -79 -91
rect -113 -125 -79 -119
rect -113 -187 -79 -163
rect -113 -197 -79 -187
rect -113 -255 -79 -235
rect -113 -269 -79 -255
rect -113 -323 -79 -307
rect -113 -341 -79 -323
rect -113 -391 -79 -379
rect -113 -413 -79 -391
rect -17 391 17 413
rect -17 379 17 391
rect -17 323 17 341
rect -17 307 17 323
rect -17 255 17 269
rect -17 235 17 255
rect -17 187 17 197
rect -17 163 17 187
rect -17 119 17 125
rect -17 91 17 119
rect -17 51 17 53
rect -17 19 17 51
rect -17 -51 17 -19
rect -17 -53 17 -51
rect -17 -119 17 -91
rect -17 -125 17 -119
rect -17 -187 17 -163
rect -17 -197 17 -187
rect -17 -255 17 -235
rect -17 -269 17 -255
rect -17 -323 17 -307
rect -17 -341 17 -323
rect -17 -391 17 -379
rect -17 -413 17 -391
rect 79 391 113 413
rect 79 379 113 391
rect 79 323 113 341
rect 79 307 113 323
rect 79 255 113 269
rect 79 235 113 255
rect 79 187 113 197
rect 79 163 113 187
rect 79 119 113 125
rect 79 91 113 119
rect 79 51 113 53
rect 79 19 113 51
rect 79 -51 113 -19
rect 79 -53 113 -51
rect 79 -119 113 -91
rect 79 -125 113 -119
rect 79 -187 113 -163
rect 79 -197 113 -187
rect 79 -255 113 -235
rect 79 -269 113 -255
rect 79 -323 113 -307
rect 79 -341 113 -323
rect 79 -391 113 -379
rect 79 -413 113 -391
<< metal1 >>
rect -119 413 -73 450
rect -119 379 -113 413
rect -79 379 -73 413
rect -119 341 -73 379
rect -119 307 -113 341
rect -79 307 -73 341
rect -119 269 -73 307
rect -119 235 -113 269
rect -79 235 -73 269
rect -119 197 -73 235
rect -119 163 -113 197
rect -79 163 -73 197
rect -119 125 -73 163
rect -119 91 -113 125
rect -79 91 -73 125
rect -119 53 -73 91
rect -119 19 -113 53
rect -79 19 -73 53
rect -119 -19 -73 19
rect -119 -53 -113 -19
rect -79 -53 -73 -19
rect -119 -91 -73 -53
rect -119 -125 -113 -91
rect -79 -125 -73 -91
rect -119 -163 -73 -125
rect -119 -197 -113 -163
rect -79 -197 -73 -163
rect -119 -235 -73 -197
rect -119 -269 -113 -235
rect -79 -269 -73 -235
rect -119 -307 -73 -269
rect -119 -341 -113 -307
rect -79 -341 -73 -307
rect -119 -379 -73 -341
rect -119 -413 -113 -379
rect -79 -413 -73 -379
rect -119 -450 -73 -413
rect -23 413 23 450
rect -23 379 -17 413
rect 17 379 23 413
rect -23 341 23 379
rect -23 307 -17 341
rect 17 307 23 341
rect -23 269 23 307
rect -23 235 -17 269
rect 17 235 23 269
rect -23 197 23 235
rect -23 163 -17 197
rect 17 163 23 197
rect -23 125 23 163
rect -23 91 -17 125
rect 17 91 23 125
rect -23 53 23 91
rect -23 19 -17 53
rect 17 19 23 53
rect -23 -19 23 19
rect -23 -53 -17 -19
rect 17 -53 23 -19
rect -23 -91 23 -53
rect -23 -125 -17 -91
rect 17 -125 23 -91
rect -23 -163 23 -125
rect -23 -197 -17 -163
rect 17 -197 23 -163
rect -23 -235 23 -197
rect -23 -269 -17 -235
rect 17 -269 23 -235
rect -23 -307 23 -269
rect -23 -341 -17 -307
rect 17 -341 23 -307
rect -23 -379 23 -341
rect -23 -413 -17 -379
rect 17 -413 23 -379
rect -23 -450 23 -413
rect 73 413 119 450
rect 73 379 79 413
rect 113 379 119 413
rect 73 341 119 379
rect 73 307 79 341
rect 113 307 119 341
rect 73 269 119 307
rect 73 235 79 269
rect 113 235 119 269
rect 73 197 119 235
rect 73 163 79 197
rect 113 163 119 197
rect 73 125 119 163
rect 73 91 79 125
rect 113 91 119 125
rect 73 53 119 91
rect 73 19 79 53
rect 113 19 119 53
rect 73 -19 119 19
rect 73 -53 79 -19
rect 113 -53 119 -19
rect 73 -91 119 -53
rect 73 -125 79 -91
rect 113 -125 119 -91
rect 73 -163 119 -125
rect 73 -197 79 -163
rect 113 -197 119 -163
rect 73 -235 119 -197
rect 73 -269 79 -235
rect 113 -269 119 -235
rect 73 -307 119 -269
rect 73 -341 79 -307
rect 113 -341 119 -307
rect 73 -379 119 -341
rect 73 -413 79 -379
rect 113 -413 119 -379
rect 73 -450 119 -413
<< end >>
