magic
tech sky130A
magscale 1 2
timestamp 1756008383
<< nwell >>
rect -36 502 182 730
rect -16 478 152 502
rect 12 444 46 478
<< pwell >>
rect -106 -254 208 -2
<< psubdiff >>
rect -80 -69 182 -28
rect -80 -103 -61 -69
rect -27 -103 31 -69
rect 65 -103 123 -69
rect 157 -103 182 -69
rect -80 -161 182 -103
rect -80 -195 -61 -161
rect -27 -195 31 -161
rect 65 -195 123 -161
rect 157 -195 182 -161
rect -80 -228 182 -195
<< nsubdiff >>
rect 0 663 146 694
rect 0 629 29 663
rect 63 629 146 663
rect 0 571 146 629
rect 0 537 29 571
rect 63 537 146 571
rect 0 494 146 537
<< psubdiffcont >>
rect -61 -103 -27 -69
rect 31 -103 65 -69
rect 123 -103 157 -69
rect -61 -195 -27 -161
rect 31 -195 65 -161
rect 123 -195 157 -161
<< nsubdiffcont >>
rect 29 629 63 663
rect 29 537 63 571
<< poly >>
rect -80 188 -14 204
rect 58 188 88 214
rect -80 187 88 188
rect -80 153 -64 187
rect -30 153 88 187
rect -80 148 88 153
rect -80 136 -14 148
rect 58 136 88 148
<< polycont >>
rect -64 153 -30 187
<< locali >>
rect -80 663 182 680
rect -80 629 -63 663
rect -29 629 29 663
rect 63 629 121 663
rect 155 629 182 663
rect -80 571 182 629
rect -80 537 -63 571
rect -29 537 29 571
rect 63 537 121 571
rect 155 537 182 571
rect -80 508 182 537
rect 12 444 46 508
rect -80 187 -14 204
rect -80 153 -64 187
rect -30 153 -14 187
rect -80 136 -14 153
rect 100 188 134 236
rect 100 148 182 188
rect 100 114 134 148
rect 12 -44 46 22
rect -80 -69 182 -44
rect -80 -103 -61 -69
rect -27 -103 31 -69
rect 65 -103 123 -69
rect 157 -103 182 -69
rect -80 -161 182 -103
rect -80 -195 -61 -161
rect -27 -195 31 -161
rect 65 -195 123 -161
rect 157 -195 182 -161
rect -80 -212 182 -195
<< viali >>
rect -63 629 -29 663
rect 29 629 63 663
rect 121 629 155 663
rect -63 537 -29 571
rect 29 537 63 571
rect 121 537 155 571
rect -61 -103 -27 -69
rect 31 -103 65 -69
rect 123 -103 157 -69
rect -61 -195 -27 -161
rect 31 -195 65 -161
rect 123 -195 157 -161
<< metal1 >>
rect -80 663 182 680
rect -80 629 -63 663
rect -29 629 29 663
rect 63 629 121 663
rect 155 629 182 663
rect -80 571 182 629
rect -80 537 -63 571
rect -29 537 29 571
rect 63 537 121 571
rect 155 537 182 571
rect -80 508 182 537
rect -80 -69 182 -44
rect -80 -103 -61 -69
rect -27 -103 31 -69
rect 65 -103 123 -69
rect 157 -103 182 -69
rect -80 -161 182 -103
rect -80 -195 -61 -161
rect -27 -195 31 -161
rect 65 -195 123 -161
rect 157 -195 182 -161
rect -80 -212 182 -195
use sky130_fd_pr__nfet_01v8_PNPQML  sky130_fd_pr__nfet_01v8_PNPQML_0
timestamp 1756008383
transform 1 0 73 0 1 68
box -99 -68 99 68
use sky130_fd_pr__pfet_01v8_TH65V5  sky130_fd_pr__pfet_01v8_TH65V5_0
timestamp 1756008383
transform 1 0 73 0 1 340
box -109 -162 109 162
<< end >>
