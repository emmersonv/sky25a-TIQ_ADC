magic
tech sky130A
magscale 1 2
timestamp 1756008383
<< nwell >>
rect 200 856 236 892
rect 278 856 314 892
rect 462 856 498 892
rect 540 856 576 892
rect 200 764 236 800
rect 278 764 314 800
rect 462 764 498 800
rect 540 764 576 800
rect 200 -128 236 -92
rect 278 -128 314 -92
rect 462 -128 498 -92
rect 540 -128 576 -92
rect 200 -220 236 -184
rect 278 -220 314 -184
rect 462 -220 498 -184
rect 540 -220 576 -184
rect 200 -1114 236 -1078
rect 278 -1114 314 -1078
rect 462 -1114 498 -1078
rect 540 -1114 576 -1078
rect 200 -1206 236 -1170
rect 278 -1206 314 -1170
rect 462 -1206 498 -1170
rect 540 -1206 576 -1170
rect 200 -2098 236 -2062
rect 278 -2098 314 -2062
rect 462 -2098 498 -2062
rect 540 -2098 576 -2062
rect 200 -2190 236 -2154
rect 278 -2190 314 -2154
rect 462 -2190 498 -2154
rect 540 -2190 576 -2154
rect 200 -3082 236 -3046
rect 278 -3082 314 -3046
rect 462 -3082 498 -3046
rect 540 -3082 576 -3046
rect 200 -3174 236 -3138
rect 278 -3174 314 -3138
rect 462 -3174 498 -3138
rect 540 -3174 576 -3138
rect 200 -4066 236 -4030
rect 278 -4066 314 -4030
rect 462 -4066 498 -4030
rect 540 -4066 576 -4030
rect 200 -4158 236 -4122
rect 278 -4158 314 -4122
rect 462 -4158 498 -4122
rect 540 -4158 576 -4122
rect 200 -5050 236 -5014
rect 278 -5050 314 -5014
rect 462 -5050 498 -5014
rect 540 -5050 576 -5014
rect 200 -5142 236 -5106
rect 278 -5142 314 -5106
rect 462 -5142 498 -5106
rect 540 -5142 576 -5106
<< pwell >>
rect -26 -10 812 210
rect -26 -994 812 -774
rect -28 -1980 814 -1758
rect -26 -2966 812 -2744
rect -26 -3948 812 -3728
rect -26 -4932 812 -4710
rect -26 -5916 812 -5696
<< psubdiff >>
rect 0 16 786 184
rect 0 -968 786 -800
rect -2 -1954 788 -1784
rect 0 -2940 786 -2770
rect 0 -3922 786 -3754
rect 0 -4906 786 -4736
rect 0 -5890 786 -5722
<< nsubdiff >>
rect 200 891 236 892
rect 200 857 201 891
rect 235 857 236 891
rect 200 856 236 857
rect 278 891 314 892
rect 278 857 279 891
rect 313 857 314 891
rect 278 856 314 857
rect 462 891 498 892
rect 462 857 463 891
rect 497 857 498 891
rect 462 856 498 857
rect 540 891 576 892
rect 540 857 541 891
rect 575 857 576 891
rect 540 856 576 857
rect 200 799 236 800
rect 200 765 201 799
rect 235 765 236 799
rect 200 764 236 765
rect 278 799 314 800
rect 278 765 279 799
rect 313 765 314 799
rect 278 764 314 765
rect 462 799 498 800
rect 462 765 463 799
rect 497 765 498 799
rect 462 764 498 765
rect 540 799 576 800
rect 540 765 541 799
rect 575 765 576 799
rect 540 764 576 765
rect 200 -93 236 -92
rect 200 -127 201 -93
rect 235 -127 236 -93
rect 200 -128 236 -127
rect 278 -93 314 -92
rect 278 -127 279 -93
rect 313 -127 314 -93
rect 278 -128 314 -127
rect 462 -93 498 -92
rect 462 -127 463 -93
rect 497 -127 498 -93
rect 462 -128 498 -127
rect 540 -93 576 -92
rect 540 -127 541 -93
rect 575 -127 576 -93
rect 540 -128 576 -127
rect 200 -185 236 -184
rect 200 -219 201 -185
rect 235 -219 236 -185
rect 200 -220 236 -219
rect 278 -185 314 -184
rect 278 -219 279 -185
rect 313 -219 314 -185
rect 278 -220 314 -219
rect 462 -185 498 -184
rect 462 -219 463 -185
rect 497 -219 498 -185
rect 462 -220 498 -219
rect 540 -185 576 -184
rect 540 -219 541 -185
rect 575 -219 576 -185
rect 540 -220 576 -219
rect 200 -1079 236 -1078
rect 200 -1113 201 -1079
rect 235 -1113 236 -1079
rect 200 -1114 236 -1113
rect 278 -1079 314 -1078
rect 278 -1113 279 -1079
rect 313 -1113 314 -1079
rect 278 -1114 314 -1113
rect 462 -1079 498 -1078
rect 462 -1113 463 -1079
rect 497 -1113 498 -1079
rect 462 -1114 498 -1113
rect 540 -1079 576 -1078
rect 540 -1113 541 -1079
rect 575 -1113 576 -1079
rect 540 -1114 576 -1113
rect 200 -1171 236 -1170
rect 200 -1205 201 -1171
rect 235 -1205 236 -1171
rect 200 -1206 236 -1205
rect 278 -1171 314 -1170
rect 278 -1205 279 -1171
rect 313 -1205 314 -1171
rect 278 -1206 314 -1205
rect 462 -1171 498 -1170
rect 462 -1205 463 -1171
rect 497 -1205 498 -1171
rect 462 -1206 498 -1205
rect 540 -1171 576 -1170
rect 540 -1205 541 -1171
rect 575 -1205 576 -1171
rect 540 -1206 576 -1205
rect 200 -2063 236 -2062
rect 200 -2097 201 -2063
rect 235 -2097 236 -2063
rect 200 -2098 236 -2097
rect 278 -2063 314 -2062
rect 278 -2097 279 -2063
rect 313 -2097 314 -2063
rect 278 -2098 314 -2097
rect 462 -2063 498 -2062
rect 462 -2097 463 -2063
rect 497 -2097 498 -2063
rect 462 -2098 498 -2097
rect 540 -2063 576 -2062
rect 540 -2097 541 -2063
rect 575 -2097 576 -2063
rect 540 -2098 576 -2097
rect 200 -2155 236 -2154
rect 200 -2189 201 -2155
rect 235 -2189 236 -2155
rect 200 -2190 236 -2189
rect 278 -2155 314 -2154
rect 278 -2189 279 -2155
rect 313 -2189 314 -2155
rect 278 -2190 314 -2189
rect 462 -2155 498 -2154
rect 462 -2189 463 -2155
rect 497 -2189 498 -2155
rect 462 -2190 498 -2189
rect 540 -2155 576 -2154
rect 540 -2189 541 -2155
rect 575 -2189 576 -2155
rect 540 -2190 576 -2189
rect 200 -3047 236 -3046
rect 200 -3081 201 -3047
rect 235 -3081 236 -3047
rect 200 -3082 236 -3081
rect 278 -3047 314 -3046
rect 278 -3081 279 -3047
rect 313 -3081 314 -3047
rect 278 -3082 314 -3081
rect 462 -3047 498 -3046
rect 462 -3081 463 -3047
rect 497 -3081 498 -3047
rect 462 -3082 498 -3081
rect 540 -3047 576 -3046
rect 540 -3081 541 -3047
rect 575 -3081 576 -3047
rect 540 -3082 576 -3081
rect 200 -3139 236 -3138
rect 200 -3173 201 -3139
rect 235 -3173 236 -3139
rect 200 -3174 236 -3173
rect 278 -3139 314 -3138
rect 278 -3173 279 -3139
rect 313 -3173 314 -3139
rect 278 -3174 314 -3173
rect 462 -3139 498 -3138
rect 462 -3173 463 -3139
rect 497 -3173 498 -3139
rect 462 -3174 498 -3173
rect 540 -3139 576 -3138
rect 540 -3173 541 -3139
rect 575 -3173 576 -3139
rect 540 -3174 576 -3173
rect 200 -4031 236 -4030
rect 200 -4065 201 -4031
rect 235 -4065 236 -4031
rect 200 -4066 236 -4065
rect 278 -4031 314 -4030
rect 278 -4065 279 -4031
rect 313 -4065 314 -4031
rect 278 -4066 314 -4065
rect 462 -4031 498 -4030
rect 462 -4065 463 -4031
rect 497 -4065 498 -4031
rect 462 -4066 498 -4065
rect 540 -4031 576 -4030
rect 540 -4065 541 -4031
rect 575 -4065 576 -4031
rect 540 -4066 576 -4065
rect 200 -4123 236 -4122
rect 200 -4157 201 -4123
rect 235 -4157 236 -4123
rect 200 -4158 236 -4157
rect 278 -4123 314 -4122
rect 278 -4157 279 -4123
rect 313 -4157 314 -4123
rect 278 -4158 314 -4157
rect 462 -4123 498 -4122
rect 462 -4157 463 -4123
rect 497 -4157 498 -4123
rect 462 -4158 498 -4157
rect 540 -4123 576 -4122
rect 540 -4157 541 -4123
rect 575 -4157 576 -4123
rect 540 -4158 576 -4157
rect 200 -5015 236 -5014
rect 200 -5049 201 -5015
rect 235 -5049 236 -5015
rect 200 -5050 236 -5049
rect 278 -5015 314 -5014
rect 278 -5049 279 -5015
rect 313 -5049 314 -5015
rect 278 -5050 314 -5049
rect 462 -5015 498 -5014
rect 462 -5049 463 -5015
rect 497 -5049 498 -5015
rect 462 -5050 498 -5049
rect 540 -5015 576 -5014
rect 540 -5049 541 -5015
rect 575 -5049 576 -5015
rect 540 -5050 576 -5049
rect 200 -5107 236 -5106
rect 200 -5141 201 -5107
rect 235 -5141 236 -5107
rect 200 -5142 236 -5141
rect 278 -5107 314 -5106
rect 278 -5141 279 -5107
rect 313 -5141 314 -5107
rect 278 -5142 314 -5141
rect 462 -5107 498 -5106
rect 462 -5141 463 -5107
rect 497 -5141 498 -5107
rect 462 -5142 498 -5141
rect 540 -5107 576 -5106
rect 540 -5141 541 -5107
rect 575 -5141 576 -5107
rect 540 -5142 576 -5141
<< nsubdiffcont >>
rect 201 857 235 891
rect 279 857 313 891
rect 463 857 497 891
rect 541 857 575 891
rect 201 765 235 799
rect 279 765 313 799
rect 463 765 497 799
rect 541 765 575 799
rect 201 -127 235 -93
rect 279 -127 313 -93
rect 463 -127 497 -93
rect 541 -127 575 -93
rect 201 -219 235 -185
rect 279 -219 313 -185
rect 463 -219 497 -185
rect 541 -219 575 -185
rect 201 -1113 235 -1079
rect 279 -1113 313 -1079
rect 463 -1113 497 -1079
rect 541 -1113 575 -1079
rect 201 -1205 235 -1171
rect 279 -1205 313 -1171
rect 463 -1205 497 -1171
rect 541 -1205 575 -1171
rect 201 -2097 235 -2063
rect 279 -2097 313 -2063
rect 463 -2097 497 -2063
rect 541 -2097 575 -2063
rect 201 -2189 235 -2155
rect 279 -2189 313 -2155
rect 463 -2189 497 -2155
rect 541 -2189 575 -2155
rect 201 -3081 235 -3047
rect 279 -3081 313 -3047
rect 463 -3081 497 -3047
rect 541 -3081 575 -3047
rect 201 -3173 235 -3139
rect 279 -3173 313 -3139
rect 463 -3173 497 -3139
rect 541 -3173 575 -3139
rect 201 -4065 235 -4031
rect 279 -4065 313 -4031
rect 463 -4065 497 -4031
rect 541 -4065 575 -4031
rect 201 -4157 235 -4123
rect 279 -4157 313 -4123
rect 463 -4157 497 -4123
rect 541 -4157 575 -4123
rect 201 -5049 235 -5015
rect 279 -5049 313 -5015
rect 463 -5049 497 -5015
rect 541 -5049 575 -5015
rect 201 -5141 235 -5107
rect 279 -5141 313 -5107
rect 463 -5141 497 -5107
rect 541 -5141 575 -5107
<< locali >>
rect 200 891 236 892
rect 200 857 201 891
rect 235 857 236 891
rect 200 856 236 857
rect 278 891 314 892
rect 278 857 279 891
rect 313 857 314 891
rect 278 856 314 857
rect 462 891 498 892
rect 462 857 463 891
rect 497 857 498 891
rect 462 856 498 857
rect 540 891 576 892
rect 540 857 541 891
rect 575 857 576 891
rect 540 856 576 857
rect 200 799 236 800
rect 200 765 201 799
rect 235 765 236 799
rect 200 764 236 765
rect 278 799 314 800
rect 278 765 279 799
rect 313 765 314 799
rect 278 764 314 765
rect 462 799 498 800
rect 462 765 463 799
rect 497 765 498 799
rect 462 764 498 765
rect 540 799 576 800
rect 540 765 541 799
rect 575 765 576 799
rect 540 764 576 765
rect 0 364 66 432
rect 738 376 786 416
rect 0 16 786 184
rect 200 -93 236 -92
rect 200 -127 201 -93
rect 235 -127 236 -93
rect 200 -128 236 -127
rect 278 -93 314 -92
rect 278 -127 279 -93
rect 313 -127 314 -93
rect 278 -128 314 -127
rect 462 -93 498 -92
rect 462 -127 463 -93
rect 497 -127 498 -93
rect 462 -128 498 -127
rect 540 -93 576 -92
rect 540 -127 541 -93
rect 575 -127 576 -93
rect 540 -128 576 -127
rect 200 -185 236 -184
rect 200 -219 201 -185
rect 235 -219 236 -185
rect 200 -220 236 -219
rect 278 -185 314 -184
rect 278 -219 279 -185
rect 313 -219 314 -185
rect 278 -220 314 -219
rect 462 -185 498 -184
rect 462 -219 463 -185
rect 497 -219 498 -185
rect 462 -220 498 -219
rect 540 -185 576 -184
rect 540 -219 541 -185
rect 575 -219 576 -185
rect 540 -220 576 -219
rect 0 -620 66 -552
rect 738 -608 786 -568
rect 0 -968 786 -800
rect 200 -1079 236 -1078
rect 200 -1113 201 -1079
rect 235 -1113 236 -1079
rect 200 -1114 236 -1113
rect 278 -1079 314 -1078
rect 278 -1113 279 -1079
rect 313 -1113 314 -1079
rect 278 -1114 314 -1113
rect 462 -1079 498 -1078
rect 462 -1113 463 -1079
rect 497 -1113 498 -1079
rect 462 -1114 498 -1113
rect 540 -1079 576 -1078
rect 540 -1113 541 -1079
rect 575 -1113 576 -1079
rect 540 -1114 576 -1113
rect 200 -1171 236 -1170
rect 200 -1205 201 -1171
rect 235 -1205 236 -1171
rect 200 -1206 236 -1205
rect 278 -1171 314 -1170
rect 278 -1205 279 -1171
rect 313 -1205 314 -1171
rect 278 -1206 314 -1205
rect 462 -1171 498 -1170
rect 462 -1205 463 -1171
rect 497 -1205 498 -1171
rect 462 -1206 498 -1205
rect 540 -1171 576 -1170
rect 540 -1205 541 -1171
rect 575 -1205 576 -1171
rect 540 -1206 576 -1205
rect 0 -1606 66 -1538
rect 738 -1594 786 -1554
rect -2 -1954 788 -1784
rect 200 -2063 236 -2062
rect 200 -2097 201 -2063
rect 235 -2097 236 -2063
rect 200 -2098 236 -2097
rect 278 -2063 314 -2062
rect 278 -2097 279 -2063
rect 313 -2097 314 -2063
rect 278 -2098 314 -2097
rect 462 -2063 498 -2062
rect 462 -2097 463 -2063
rect 497 -2097 498 -2063
rect 462 -2098 498 -2097
rect 540 -2063 576 -2062
rect 540 -2097 541 -2063
rect 575 -2097 576 -2063
rect 540 -2098 576 -2097
rect 200 -2155 236 -2154
rect 200 -2189 201 -2155
rect 235 -2189 236 -2155
rect 200 -2190 236 -2189
rect 278 -2155 314 -2154
rect 278 -2189 279 -2155
rect 313 -2189 314 -2155
rect 278 -2190 314 -2189
rect 462 -2155 498 -2154
rect 462 -2189 463 -2155
rect 497 -2189 498 -2155
rect 462 -2190 498 -2189
rect 540 -2155 576 -2154
rect 540 -2189 541 -2155
rect 575 -2189 576 -2155
rect 540 -2190 576 -2189
rect 0 -2590 66 -2522
rect 738 -2578 786 -2538
rect 0 -2940 786 -2770
rect 200 -3047 236 -3046
rect 200 -3081 201 -3047
rect 235 -3081 236 -3047
rect 200 -3082 236 -3081
rect 278 -3047 314 -3046
rect 278 -3081 279 -3047
rect 313 -3081 314 -3047
rect 278 -3082 314 -3081
rect 462 -3047 498 -3046
rect 462 -3081 463 -3047
rect 497 -3081 498 -3047
rect 462 -3082 498 -3081
rect 540 -3047 576 -3046
rect 540 -3081 541 -3047
rect 575 -3081 576 -3047
rect 540 -3082 576 -3081
rect 200 -3139 236 -3138
rect 200 -3173 201 -3139
rect 235 -3173 236 -3139
rect 200 -3174 236 -3173
rect 278 -3139 314 -3138
rect 278 -3173 279 -3139
rect 313 -3173 314 -3139
rect 278 -3174 314 -3173
rect 462 -3139 498 -3138
rect 462 -3173 463 -3139
rect 497 -3173 498 -3139
rect 462 -3174 498 -3173
rect 540 -3139 576 -3138
rect 540 -3173 541 -3139
rect 575 -3173 576 -3139
rect 540 -3174 576 -3173
rect 0 -3574 66 -3506
rect 738 -3562 786 -3522
rect 0 -3922 786 -3754
rect 200 -4031 236 -4030
rect 200 -4065 201 -4031
rect 235 -4065 236 -4031
rect 200 -4066 236 -4065
rect 278 -4031 314 -4030
rect 278 -4065 279 -4031
rect 313 -4065 314 -4031
rect 278 -4066 314 -4065
rect 462 -4031 498 -4030
rect 462 -4065 463 -4031
rect 497 -4065 498 -4031
rect 462 -4066 498 -4065
rect 540 -4031 576 -4030
rect 540 -4065 541 -4031
rect 575 -4065 576 -4031
rect 540 -4066 576 -4065
rect 200 -4123 236 -4122
rect 200 -4157 201 -4123
rect 235 -4157 236 -4123
rect 200 -4158 236 -4157
rect 278 -4123 314 -4122
rect 278 -4157 279 -4123
rect 313 -4157 314 -4123
rect 278 -4158 314 -4157
rect 462 -4123 498 -4122
rect 462 -4157 463 -4123
rect 497 -4157 498 -4123
rect 462 -4158 498 -4157
rect 540 -4123 576 -4122
rect 540 -4157 541 -4123
rect 575 -4157 576 -4123
rect 540 -4158 576 -4157
rect 0 -4558 66 -4490
rect 738 -4546 786 -4506
rect 0 -4906 786 -4736
rect 200 -5015 236 -5014
rect 200 -5049 201 -5015
rect 235 -5049 236 -5015
rect 200 -5050 236 -5049
rect 278 -5015 314 -5014
rect 278 -5049 279 -5015
rect 313 -5049 314 -5015
rect 278 -5050 314 -5049
rect 462 -5015 498 -5014
rect 462 -5049 463 -5015
rect 497 -5049 498 -5015
rect 462 -5050 498 -5049
rect 540 -5015 576 -5014
rect 540 -5049 541 -5015
rect 575 -5049 576 -5015
rect 540 -5050 576 -5049
rect 200 -5107 236 -5106
rect 200 -5141 201 -5107
rect 235 -5141 236 -5107
rect 200 -5142 236 -5141
rect 278 -5107 314 -5106
rect 278 -5141 279 -5107
rect 313 -5141 314 -5107
rect 278 -5142 314 -5141
rect 462 -5107 498 -5106
rect 462 -5141 463 -5107
rect 497 -5141 498 -5107
rect 462 -5142 498 -5141
rect 540 -5107 576 -5106
rect 540 -5141 541 -5107
rect 575 -5141 576 -5107
rect 540 -5142 576 -5141
rect 0 -5542 66 -5474
rect 738 -5530 786 -5490
rect 0 -5890 786 -5722
<< viali >>
rect 201 857 235 891
rect 279 857 313 891
rect 463 857 497 891
rect 541 857 575 891
rect 201 765 235 799
rect 279 765 313 799
rect 463 765 497 799
rect 541 765 575 799
rect 201 -127 235 -93
rect 279 -127 313 -93
rect 463 -127 497 -93
rect 541 -127 575 -93
rect 201 -219 235 -185
rect 279 -219 313 -185
rect 463 -219 497 -185
rect 541 -219 575 -185
rect 201 -1113 235 -1079
rect 279 -1113 313 -1079
rect 463 -1113 497 -1079
rect 541 -1113 575 -1079
rect 201 -1205 235 -1171
rect 279 -1205 313 -1171
rect 463 -1205 497 -1171
rect 541 -1205 575 -1171
rect 201 -2097 235 -2063
rect 279 -2097 313 -2063
rect 463 -2097 497 -2063
rect 541 -2097 575 -2063
rect 201 -2189 235 -2155
rect 279 -2189 313 -2155
rect 463 -2189 497 -2155
rect 541 -2189 575 -2155
rect 201 -3081 235 -3047
rect 279 -3081 313 -3047
rect 463 -3081 497 -3047
rect 541 -3081 575 -3047
rect 201 -3173 235 -3139
rect 279 -3173 313 -3139
rect 463 -3173 497 -3139
rect 541 -3173 575 -3139
rect 201 -4065 235 -4031
rect 279 -4065 313 -4031
rect 463 -4065 497 -4031
rect 541 -4065 575 -4031
rect 201 -4157 235 -4123
rect 279 -4157 313 -4123
rect 463 -4157 497 -4123
rect 541 -4157 575 -4123
rect 201 -5049 235 -5015
rect 279 -5049 313 -5015
rect 463 -5049 497 -5015
rect 541 -5049 575 -5015
rect 201 -5141 235 -5107
rect 279 -5141 313 -5107
rect 463 -5141 497 -5107
rect 541 -5141 575 -5107
<< metal1 >>
rect 0 891 788 908
rect 0 857 201 891
rect 235 857 279 891
rect 313 857 463 891
rect 497 857 541 891
rect 575 857 788 891
rect 0 799 788 857
rect 0 765 201 799
rect 235 765 279 799
rect 313 765 463 799
rect 497 765 541 799
rect 575 765 788 799
rect 0 736 788 765
rect 0 16 786 184
rect 2 -93 790 -74
rect 2 -127 201 -93
rect 235 -127 279 -93
rect 313 -127 463 -93
rect 497 -127 541 -93
rect 575 -127 790 -93
rect 2 -185 790 -127
rect 2 -219 201 -185
rect 235 -219 279 -185
rect 313 -219 463 -185
rect 497 -219 541 -185
rect 575 -219 790 -185
rect 2 -246 790 -219
rect 0 -968 786 -800
rect 0 -1079 788 -1062
rect 0 -1113 201 -1079
rect 235 -1113 279 -1079
rect 313 -1113 463 -1079
rect 497 -1113 541 -1079
rect 575 -1113 788 -1079
rect 0 -1171 788 -1113
rect 0 -1205 201 -1171
rect 235 -1205 279 -1171
rect 313 -1205 463 -1171
rect 497 -1205 541 -1171
rect 575 -1205 788 -1171
rect 0 -1234 788 -1205
rect -2 -1954 788 -1784
rect 0 -2063 788 -2046
rect 0 -2097 201 -2063
rect 235 -2097 279 -2063
rect 313 -2097 463 -2063
rect 497 -2097 541 -2063
rect 575 -2097 788 -2063
rect 0 -2155 788 -2097
rect 0 -2189 201 -2155
rect 235 -2189 279 -2155
rect 313 -2189 463 -2155
rect 497 -2189 541 -2155
rect 575 -2189 788 -2155
rect 0 -2218 788 -2189
rect 0 -2940 786 -2770
rect 0 -3047 788 -3030
rect 0 -3081 201 -3047
rect 235 -3081 279 -3047
rect 313 -3081 463 -3047
rect 497 -3081 541 -3047
rect 575 -3081 788 -3047
rect 0 -3139 788 -3081
rect 0 -3173 201 -3139
rect 235 -3173 279 -3139
rect 313 -3173 463 -3139
rect 497 -3173 541 -3139
rect 575 -3173 788 -3139
rect 0 -3202 788 -3173
rect 0 -3922 786 -3754
rect 0 -4031 788 -4014
rect 0 -4065 201 -4031
rect 235 -4065 279 -4031
rect 313 -4065 463 -4031
rect 497 -4065 541 -4031
rect 575 -4065 788 -4031
rect 0 -4123 788 -4065
rect 0 -4157 201 -4123
rect 235 -4157 279 -4123
rect 313 -4157 463 -4123
rect 497 -4157 541 -4123
rect 575 -4157 788 -4123
rect 0 -4186 788 -4157
rect 0 -4906 786 -4736
rect 0 -5015 788 -4998
rect 0 -5049 201 -5015
rect 235 -5049 279 -5015
rect 313 -5049 463 -5015
rect 497 -5049 541 -5015
rect 575 -5049 788 -5015
rect 0 -5107 788 -5049
rect 0 -5141 201 -5107
rect 235 -5141 279 -5107
rect 313 -5141 463 -5107
rect 497 -5141 541 -5107
rect 575 -5141 788 -5107
rect 0 -5170 788 -5141
rect 0 -5890 786 -5722
use gain_stage  gain_stage_0
timestamp 1756008383
transform 1 0 0 0 1 0
box -26 -26 812 958
use gain_stage  gain_stage_1
timestamp 1756008383
transform 1 0 0 0 1 -984
box -26 -26 812 958
use gain_stage  gain_stage_2
timestamp 1756008383
transform 1 0 0 0 1 -1970
box -26 -26 812 958
use gain_stage  gain_stage_3
timestamp 1756008383
transform 1 0 0 0 1 -2954
box -26 -26 812 958
use gain_stage  gain_stage_4
timestamp 1756008383
transform 1 0 0 0 1 -3938
box -26 -26 812 958
use gain_stage  gain_stage_5
timestamp 1756008383
transform 1 0 0 0 1 -4922
box -26 -26 812 958
use gain_stage  gain_stage_6
timestamp 1756008383
transform 1 0 0 0 1 -5906
box -26 -26 812 958
<< end >>
