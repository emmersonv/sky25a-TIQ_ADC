** sch_path: /foss/designs/analog-circuit-design/sky25a-TIQ_ADC/xschem/INVERTER_SIZES/inverter_p12_n3_symsch.sch
.subckt inverter_p12_n3_symsch Vout Vin VDPWR VGND
*.PININFO Vout:O Vin:I VDPWR:B VGND:B
x1 VDPWR Vout Vin VGND inverter_p12_n3
.ends

* expanding   symbol:  /foss/designs/analog-circuit-design/sky25a-TIQ_ADC/xschem/INVERTER_SIZES/inverter_p12_n3.sym # of pins=4
** sym_path: /foss/designs/analog-circuit-design/sky25a-TIQ_ADC/xschem/INVERTER_SIZES/inverter_p12_n3.sym
** sch_path: /foss/designs/analog-circuit-design/sky25a-TIQ_ADC/xschem/INVERTER_SIZES/inverter_p12_n3.sch
.subckt inverter_p12_n3 VDPWR Vout Vin VGND
*.PININFO Vout:O Vin:I VDPWR:B VGND:B
XM1 Vout Vin VGND VGND sky130_fd_pr__nfet_01v8 L=0.15 W=3 nf=1 m=1
XM2 Vout Vin VDPWR VDPWR sky130_fd_pr__pfet_01v8 L=0.15 W=12 nf=2 m=1
.ends

