magic
tech sky130A
magscale 1 2
timestamp 1754164428
<< nwell >>
rect -36 1490 894 3830
<< psubdiff >>
rect -36 2 894 34
rect -36 -34 30 2
rect 66 -34 122 2
rect 158 -34 214 2
rect 250 -34 306 2
rect 342 -34 398 2
rect 434 -34 490 2
rect 526 -34 582 2
rect 618 -34 674 2
rect 710 -34 766 2
rect 802 -34 894 2
rect -36 -90 894 -34
rect -36 -126 30 -90
rect 66 -126 122 -90
rect 158 -126 214 -90
rect 250 -126 306 -90
rect 342 -126 398 -90
rect 434 -126 490 -90
rect 526 -126 582 -90
rect 618 -126 674 -90
rect 710 -126 766 -90
rect 802 -126 894 -90
rect -36 -166 894 -126
<< nsubdiff >>
rect 0 3764 858 3794
rect 0 3728 64 3764
rect 100 3728 156 3764
rect 192 3728 248 3764
rect 284 3728 340 3764
rect 376 3728 432 3764
rect 468 3728 524 3764
rect 560 3728 616 3764
rect 652 3728 708 3764
rect 744 3728 800 3764
rect 836 3728 858 3764
rect 0 3672 858 3728
rect 0 3636 64 3672
rect 100 3636 156 3672
rect 192 3636 248 3672
rect 284 3636 340 3672
rect 376 3636 432 3672
rect 468 3636 524 3672
rect 560 3636 616 3672
rect 652 3636 708 3672
rect 744 3636 800 3672
rect 836 3636 858 3672
rect 0 3594 858 3636
<< psubdiffcont >>
rect 30 -34 66 2
rect 122 -34 158 2
rect 214 -34 250 2
rect 306 -34 342 2
rect 398 -34 434 2
rect 490 -34 526 2
rect 582 -34 618 2
rect 674 -34 710 2
rect 766 -34 802 2
rect 30 -126 66 -90
rect 122 -126 158 -90
rect 214 -126 250 -90
rect 306 -126 342 -90
rect 398 -126 434 -90
rect 490 -126 526 -90
rect 582 -126 618 -90
rect 674 -126 710 -90
rect 766 -126 802 -90
<< nsubdiffcont >>
rect 64 3728 100 3764
rect 156 3728 192 3764
rect 248 3728 284 3764
rect 340 3728 376 3764
rect 432 3728 468 3764
rect 524 3728 560 3764
rect 616 3728 652 3764
rect 708 3728 744 3764
rect 800 3728 836 3764
rect 64 3636 100 3672
rect 156 3636 192 3672
rect 248 3636 284 3672
rect 340 3636 376 3672
rect 432 3636 468 3672
rect 524 3636 560 3672
rect 616 3636 652 3672
rect 708 3636 744 3672
rect 800 3636 836 3672
<< poly >>
rect 0 1510 66 1526
rect 0 1476 16 1510
rect 50 1490 66 1510
rect 370 1490 400 1526
rect 50 1476 796 1490
rect 0 1460 796 1476
rect 188 1448 366 1460
rect 492 1448 670 1460
<< polycont >>
rect 16 1476 50 1510
<< locali >>
rect -36 3764 894 3780
rect -36 3728 64 3764
rect 100 3728 156 3764
rect 192 3728 248 3764
rect 284 3728 340 3764
rect 376 3728 432 3764
rect 468 3728 524 3764
rect 560 3728 616 3764
rect 652 3728 708 3764
rect 744 3728 800 3764
rect 836 3728 894 3764
rect -36 3672 894 3728
rect -36 3636 64 3672
rect 100 3636 156 3672
rect 192 3636 248 3672
rect 284 3636 340 3672
rect 376 3636 432 3672
rect 468 3636 524 3672
rect 560 3636 616 3672
rect 652 3636 708 3672
rect 744 3636 800 3672
rect 836 3636 894 3672
rect -36 3608 894 3636
rect 324 1650 358 3608
rect 0 1510 66 1526
rect 0 1476 16 1510
rect 50 1476 66 1510
rect 412 1500 446 1548
rect 792 1510 858 1526
rect 792 1500 808 1510
rect 0 1460 66 1476
rect 108 1476 808 1500
rect 842 1476 858 1510
rect 108 1460 858 1476
rect 108 1426 142 1460
rect 412 1426 446 1460
rect 716 1426 750 1460
rect 12 18 46 84
rect 204 18 238 84
rect 316 18 350 84
rect 508 18 542 84
rect 620 18 654 84
rect 812 18 846 84
rect -36 2 894 18
rect -36 -34 30 2
rect 66 -34 122 2
rect 158 -34 214 2
rect 250 -34 306 2
rect 342 -34 398 2
rect 434 -34 490 2
rect 526 -34 582 2
rect 618 -34 674 2
rect 710 -34 766 2
rect 802 -34 894 2
rect -36 -90 894 -34
rect -36 -126 30 -90
rect 66 -126 122 -90
rect 158 -126 214 -90
rect 250 -126 306 -90
rect 342 -126 398 -90
rect 434 -126 490 -90
rect 526 -126 582 -90
rect 618 -126 674 -90
rect 710 -126 766 -90
rect 802 -126 894 -90
rect -36 -150 894 -126
<< viali >>
rect 64 3728 100 3764
rect 156 3728 192 3764
rect 248 3728 284 3764
rect 340 3728 376 3764
rect 432 3728 468 3764
rect 524 3728 560 3764
rect 616 3728 652 3764
rect 708 3728 744 3764
rect 800 3728 836 3764
rect 64 3636 100 3672
rect 156 3636 192 3672
rect 248 3636 284 3672
rect 340 3636 376 3672
rect 432 3636 468 3672
rect 524 3636 560 3672
rect 616 3636 652 3672
rect 708 3636 744 3672
rect 800 3636 836 3672
rect 16 1476 50 1510
rect 808 1476 842 1510
rect 30 -34 66 2
rect 122 -34 158 2
rect 214 -34 250 2
rect 306 -34 342 2
rect 398 -34 434 2
rect 490 -34 526 2
rect 582 -34 618 2
rect 674 -34 710 2
rect 766 -34 802 2
rect 30 -126 66 -90
rect 122 -126 158 -90
rect 214 -126 250 -90
rect 306 -126 342 -90
rect 398 -126 434 -90
rect 490 -126 526 -90
rect 582 -126 618 -90
rect 674 -126 710 -90
rect 766 -126 802 -90
<< metal1 >>
rect -36 3764 894 3780
rect -36 3728 64 3764
rect 100 3728 156 3764
rect 192 3728 248 3764
rect 284 3728 340 3764
rect 376 3728 432 3764
rect 468 3728 524 3764
rect 560 3728 616 3764
rect 652 3728 708 3764
rect 744 3728 800 3764
rect 836 3728 894 3764
rect -36 3672 894 3728
rect -36 3636 64 3672
rect 100 3636 156 3672
rect 192 3636 248 3672
rect 284 3636 340 3672
rect 376 3636 432 3672
rect 468 3636 524 3672
rect 560 3636 616 3672
rect 652 3636 708 3672
rect 744 3636 800 3672
rect 836 3636 894 3672
rect -36 3608 894 3636
rect 0 1510 66 1526
rect 0 1476 16 1510
rect 50 1476 66 1510
rect 0 1460 66 1476
rect 792 1510 858 1526
rect 792 1476 808 1510
rect 842 1476 858 1510
rect 792 1460 858 1476
rect -36 2 894 18
rect -36 -34 30 2
rect 66 -34 122 2
rect 158 -34 214 2
rect 250 -34 306 2
rect 342 -34 398 2
rect 434 -34 490 2
rect 526 -34 582 2
rect 618 -34 674 2
rect 710 -34 766 2
rect 802 -34 894 2
rect -36 -90 894 -34
rect -36 -126 30 -90
rect 66 -126 122 -90
rect 158 -126 214 -90
rect 250 -126 306 -90
rect 342 -126 398 -90
rect 434 -126 490 -90
rect 526 -126 582 -90
rect 618 -126 674 -90
rect 710 -126 766 -90
rect 802 -126 894 -90
rect -36 -150 894 -126
use sky130_fd_pr__nfet_01v8_CTSNWR  sky130_fd_pr__nfet_01v8_CTSNWR_0
timestamp 1753585664
transform 1 0 125 0 1 755
box -125 -693 125 723
use sky130_fd_pr__nfet_01v8_CTSNWR  sky130_fd_pr__nfet_01v8_CTSNWR_1
timestamp 1753585664
transform 1 0 429 0 1 755
box -125 -693 125 723
use sky130_fd_pr__nfet_01v8_CTSNWR  sky130_fd_pr__nfet_01v8_CTSNWR_2
timestamp 1753585664
transform 1 0 733 0 1 755
box -125 -693 125 723
use sky130_fd_pr__pfet_01v8_FCTDLW  sky130_fd_pr__pfet_01v8_FCTDLW_0
timestamp 1753585664
transform 1 0 385 0 1 1599
box -109 -109 109 109
<< end >>
