magic
tech sky130A
magscale 1 2
timestamp 1752981230
<< nwell >>
rect -36 1624 896 2124
<< psubdiff >>
rect -36 2 896 34
rect -36 -134 32 2
rect 828 -134 896 2
rect -36 -166 896 -134
<< nsubdiff >>
rect 0 2008 860 2040
rect 0 1874 32 2008
rect 828 1874 860 2008
rect 0 1840 860 1874
<< psubdiffcont >>
rect 32 -134 828 2
<< nsubdiffcont >>
rect 32 1874 828 2008
<< poly >>
rect 8 1650 74 1666
rect 8 1616 24 1650
rect 58 1630 74 1650
rect 370 1630 400 1660
rect 58 1616 796 1630
rect 8 1612 796 1616
rect 8 1600 92 1612
rect 188 1582 670 1612
<< polycont >>
rect 24 1616 58 1650
<< locali >>
rect 12 2008 848 2028
rect 12 1872 32 2008
rect 828 1872 848 2008
rect 12 1852 848 1872
rect 324 1790 358 1852
rect 8 1650 74 1666
rect 8 1616 24 1650
rect 58 1616 74 1650
rect 412 1634 446 1682
rect 830 1650 896 1666
rect 830 1634 846 1650
rect 8 1600 74 1616
rect 108 1616 846 1634
rect 880 1616 896 1650
rect 108 1600 896 1616
rect 108 1594 750 1600
rect 108 1560 142 1594
rect 412 1560 446 1594
rect 716 1560 750 1594
rect 12 22 46 84
rect 204 22 238 86
rect 316 22 350 84
rect 508 22 542 84
rect 620 22 654 84
rect 812 22 846 86
rect 12 2 848 22
rect 12 -134 32 2
rect 828 -134 848 2
rect 12 -154 848 -134
<< viali >>
rect 32 1874 828 2008
rect 32 1872 828 1874
rect 24 1616 58 1650
rect 846 1616 880 1650
rect 32 -134 828 2
<< metal1 >>
rect 2 2008 860 2026
rect 2 1872 32 2008
rect 828 1872 860 2008
rect 2 1854 860 1872
rect -36 1650 74 1666
rect -36 1616 24 1650
rect 58 1616 74 1650
rect -36 1600 74 1616
rect 830 1650 896 1666
rect 830 1616 846 1650
rect 880 1616 896 1650
rect 830 1600 896 1616
rect -36 2 896 22
rect -36 -134 32 2
rect 828 -134 896 2
rect -36 -154 896 -134
use sky130_fd_pr__nfet_01v8_3LP5BP  sky130_fd_pr__nfet_01v8_3LP5BP_0
timestamp 1752972803
transform 1 0 125 0 1 822
box -125 -760 125 790
use sky130_fd_pr__nfet_01v8_3LP5BP  sky130_fd_pr__nfet_01v8_3LP5BP_1
timestamp 1752972803
transform 1 0 429 0 1 822
box -125 -760 125 790
use sky130_fd_pr__nfet_01v8_3LP5BP  sky130_fd_pr__nfet_01v8_3LP5BP_2
timestamp 1752972803
transform 1 0 733 0 1 822
box -125 -760 125 790
use sky130_fd_pr__pfet_01v8_7SLTNL  sky130_fd_pr__pfet_01v8_7SLTNL_0
timestamp 1752972140
transform 1 0 385 0 1 1736
box -109 -112 109 112
<< labels >>
rlabel metal1 8 1600 22 1614 7 Vin
port 3 w
rlabel metal1 390 1886 440 1940 1 VDPWR
port 1 n
rlabel metal1 882 1600 896 1614 3 Vout
port 2 e
rlabel metal1 392 -154 424 -122 5 VGND
port 4 s
<< end >>
