magic
tech sky130A
magscale 1 2
timestamp 1756008383
<< error_s >>
rect 3760 3540 3960 3698
rect 3996 3540 4128 3708
rect 3760 3504 4128 3540
rect 3960 3480 4128 3504
rect 3760 3444 4128 3480
rect 3760 3408 3960 3444
<< nwell >>
rect 1722 5016 1756 5036
rect 3760 4210 3960 4230
rect 2234 3602 3996 4210
rect 3760 3566 3960 3602
rect 3802 3016 3838 3052
rect 3894 3016 3930 3052
rect 1722 2564 1756 2928
rect 3760 2898 3960 3012
rect 3760 2564 3960 2646
rect 1656 2486 3996 2564
rect 3760 2450 3960 2486
rect 3760 2164 3960 2200
rect 1644 2034 3996 2164
rect 3760 1998 3960 2034
rect 3760 1408 3960 1444
rect 1644 1270 3996 1408
rect 3760 1234 3960 1270
<< pwell >>
rect -26 4148 226 4218
rect 14 4128 194 4148
rect -26 3540 226 3610
rect -26 2954 226 3038
rect 14 2932 194 2954
rect -26 2504 226 2590
rect 14 2472 194 2504
rect -26 2060 226 2146
<< psubdiff >>
rect 0 4189 200 4192
rect 0 4174 41 4189
rect 40 4155 41 4174
rect 75 4174 133 4189
rect 75 4155 76 4174
rect 40 4154 76 4155
rect 132 4155 133 4174
rect 167 4174 200 4189
rect 167 4155 168 4174
rect 132 4154 168 4155
rect 0 3566 200 3584
rect 0 2993 200 3012
rect 0 2980 41 2993
rect 40 2959 41 2980
rect 75 2980 133 2993
rect 75 2959 76 2980
rect 40 2958 76 2959
rect 132 2959 133 2980
rect 167 2980 200 2993
rect 167 2959 168 2980
rect 132 2958 168 2959
rect 0 2533 200 2564
rect 0 2530 41 2533
rect 40 2499 41 2530
rect 75 2530 133 2533
rect 75 2499 76 2530
rect 40 2498 76 2499
rect 132 2499 133 2530
rect 167 2530 200 2533
rect 167 2499 168 2530
rect 132 2498 168 2499
rect 0 2086 200 2120
<< nsubdiff >>
rect 3760 4174 3960 4230
rect 3760 3603 3960 3620
rect 3760 3569 3803 3603
rect 3837 3569 3895 3603
rect 3929 3569 3960 3603
rect 3760 3566 3960 3569
rect 3802 3051 3838 3052
rect 3802 3017 3803 3051
rect 3837 3017 3838 3051
rect 3802 3016 3838 3017
rect 3894 3051 3930 3052
rect 3894 3017 3895 3051
rect 3929 3017 3930 3051
rect 3894 3016 3930 3017
rect 3760 2959 3960 3012
rect 3760 2925 3803 2959
rect 3837 2925 3895 2959
rect 3929 2925 3960 2959
rect 3760 2898 3960 2925
rect 3802 2683 3838 2684
rect 3802 2649 3803 2683
rect 3837 2649 3838 2683
rect 3802 2648 3838 2649
rect 3894 2683 3930 2684
rect 3894 2649 3895 2683
rect 3929 2649 3930 2683
rect 3894 2648 3930 2649
rect 3760 2591 3960 2646
rect 3760 2557 3803 2591
rect 3837 2557 3895 2591
rect 3929 2557 3960 2591
rect 3760 2499 3960 2557
rect 3760 2465 3803 2499
rect 3837 2465 3895 2499
rect 3929 2465 3960 2499
rect 3760 2450 3960 2465
rect 3802 2223 3838 2224
rect 3802 2200 3803 2223
rect 3760 2189 3803 2200
rect 3837 2200 3838 2223
rect 3894 2223 3930 2224
rect 3894 2200 3895 2223
rect 3837 2189 3895 2200
rect 3929 2200 3930 2223
rect 3929 2189 3960 2200
rect 3760 2131 3960 2189
rect 3760 2097 3803 2131
rect 3837 2097 3895 2131
rect 3929 2097 3960 2131
rect 3760 2039 3960 2097
rect 3760 2005 3803 2039
rect 3837 2005 3895 2039
rect 3929 2005 3960 2039
rect 3760 1998 3960 2005
rect 3760 1395 3960 1444
rect 3760 1361 3803 1395
rect 3837 1361 3895 1395
rect 3929 1361 3960 1395
rect 3760 1303 3960 1361
rect 3760 1269 3803 1303
rect 3837 1269 3895 1303
rect 3929 1269 3960 1303
rect 3760 1234 3960 1269
<< psubdiffcont >>
rect 41 4155 75 4189
rect 133 4155 167 4189
rect 41 2959 75 2993
rect 133 2959 167 2993
rect 41 2499 75 2533
rect 133 2499 167 2533
<< nsubdiffcont >>
rect 3803 3569 3837 3603
rect 3895 3569 3929 3603
rect 3803 3017 3837 3051
rect 3895 3017 3929 3051
rect 3803 2925 3837 2959
rect 3895 2925 3929 2959
rect 3803 2649 3837 2683
rect 3895 2649 3929 2683
rect 3803 2557 3837 2591
rect 3895 2557 3929 2591
rect 3803 2465 3837 2499
rect 3895 2465 3929 2499
rect 3803 2189 3837 2223
rect 3895 2189 3929 2223
rect 3803 2097 3837 2131
rect 3895 2097 3929 2131
rect 3803 2005 3837 2039
rect 3895 2005 3929 2039
rect 3803 1361 3837 1395
rect 3895 1361 3929 1395
rect 3803 1269 3837 1303
rect 3895 1269 3929 1303
<< locali >>
rect 16 4189 184 4192
rect 16 4174 41 4189
rect 40 4155 41 4174
rect 75 4174 133 4189
rect 75 4155 76 4174
rect 40 4154 76 4155
rect 132 4155 133 4174
rect 167 4174 184 4189
rect 167 4155 168 4174
rect 132 4154 168 4155
rect 3802 3603 3838 3604
rect 3802 3569 3803 3603
rect 3837 3569 3838 3603
rect 3802 3568 3838 3569
rect 3894 3603 3930 3604
rect 3894 3569 3895 3603
rect 3929 3569 3930 3603
rect 3894 3568 3930 3569
rect 3802 3051 3838 3052
rect 3802 3017 3803 3051
rect 3837 3017 3838 3051
rect 3802 3016 3838 3017
rect 3894 3051 3930 3052
rect 3894 3017 3895 3051
rect 3929 3017 3930 3051
rect 3894 3016 3930 3017
rect 40 2993 76 2994
rect 40 2959 41 2993
rect 75 2959 76 2993
rect 40 2958 76 2959
rect 132 2993 168 2994
rect 132 2959 133 2993
rect 167 2959 168 2993
rect 132 2958 168 2959
rect 3802 2959 3838 2960
rect 3802 2925 3803 2959
rect 3837 2925 3838 2959
rect 3802 2924 3838 2925
rect 3894 2959 3930 2960
rect 3894 2925 3895 2959
rect 3929 2925 3930 2959
rect 3894 2924 3930 2925
rect 3802 2683 3838 2684
rect 3802 2649 3803 2683
rect 3837 2649 3838 2683
rect 3802 2648 3838 2649
rect 3894 2683 3930 2684
rect 3894 2649 3895 2683
rect 3929 2649 3930 2683
rect 3894 2648 3930 2649
rect 3802 2591 3838 2592
rect 3802 2564 3803 2591
rect 16 2533 184 2564
rect 16 2530 41 2533
rect 40 2499 41 2530
rect 75 2530 133 2533
rect 75 2499 76 2530
rect 40 2498 76 2499
rect 132 2499 133 2530
rect 167 2530 184 2533
rect 3774 2557 3803 2564
rect 3837 2564 3838 2591
rect 3894 2591 3930 2592
rect 3894 2564 3895 2591
rect 3837 2557 3895 2564
rect 3929 2564 3930 2591
rect 3929 2557 3946 2564
rect 167 2499 168 2530
rect 132 2498 168 2499
rect 3774 2499 3946 2557
rect 3774 2486 3803 2499
rect 3802 2465 3803 2486
rect 3837 2486 3895 2499
rect 3837 2465 3838 2486
rect 3802 2464 3838 2465
rect 3894 2465 3895 2486
rect 3929 2486 3946 2499
rect 3929 2465 3930 2486
rect 3894 2464 3930 2465
rect 3802 2223 3838 2224
rect 3802 2189 3803 2223
rect 3837 2189 3838 2223
rect 3802 2188 3838 2189
rect 3894 2223 3930 2224
rect 3894 2189 3895 2223
rect 3929 2189 3930 2223
rect 3894 2188 3930 2189
rect 3774 2131 3946 2164
rect 16 2086 184 2120
rect 3774 2097 3803 2131
rect 3837 2097 3895 2131
rect 3929 2097 3946 2131
rect 3774 2086 3946 2097
rect 3802 2039 3838 2040
rect 3802 2005 3803 2039
rect 3837 2005 3838 2039
rect 3802 2004 3838 2005
rect 3894 2039 3930 2040
rect 3894 2005 3895 2039
rect 3929 2005 3930 2039
rect 3894 2004 3930 2005
rect 3802 1395 3838 1396
rect 3802 1361 3803 1395
rect 3837 1361 3838 1395
rect 3802 1360 3838 1361
rect 3894 1395 3930 1396
rect 3894 1361 3895 1395
rect 3929 1361 3930 1395
rect 3894 1360 3930 1361
rect 3802 1303 3838 1304
rect 3802 1269 3803 1303
rect 3837 1269 3838 1303
rect 3802 1268 3838 1269
rect 3894 1303 3930 1304
rect 3894 1269 3895 1303
rect 3929 1269 3930 1303
rect 3894 1268 3930 1269
<< viali >>
rect 41 4155 75 4189
rect 133 4155 167 4189
rect 3803 3569 3837 3603
rect 3895 3569 3929 3603
rect 3803 3017 3837 3051
rect 3895 3017 3929 3051
rect 41 2959 75 2993
rect 133 2959 167 2993
rect 3803 2925 3837 2959
rect 3895 2925 3929 2959
rect 41 2499 75 2533
rect 133 2499 167 2533
rect 3803 2557 3837 2591
rect 3895 2557 3929 2591
rect 3803 2465 3837 2499
rect 3895 2465 3929 2499
rect 3803 2097 3837 2131
rect 3895 2097 3929 2131
rect 3803 1361 3837 1395
rect 3895 1361 3929 1395
rect 3803 1269 3837 1303
<< metal1 >>
rect 1632 5079 1686 5080
rect 1632 5027 1633 5079
rect 1685 5027 1686 5079
rect 1632 5026 1686 5027
rect 1632 4287 1686 4288
rect 1632 4235 1633 4287
rect 1685 4235 1686 4287
rect 1632 4234 1686 4235
rect 16 4189 184 4192
rect 16 4174 41 4189
rect 40 4155 41 4174
rect 75 4174 133 4189
rect 75 4155 76 4174
rect 40 4154 76 4155
rect 132 4155 133 4174
rect 167 4174 184 4189
rect 167 4155 168 4174
rect 132 4154 168 4155
rect 1632 4167 1686 4168
rect 1632 4115 1633 4167
rect 1685 4115 1686 4167
rect 1632 4114 1686 4115
rect 1632 3679 1686 3680
rect 1632 3627 1633 3679
rect 1685 3627 1686 3679
rect 1632 3626 1686 3627
rect 3802 3603 3838 3604
rect 3802 3569 3803 3603
rect 3837 3569 3838 3603
rect 3802 3568 3838 3569
rect 3894 3603 3930 3604
rect 3894 3569 3895 3603
rect 3929 3569 3930 3603
rect 3894 3568 3930 3569
rect 1632 3559 1686 3560
rect 1632 3507 1633 3559
rect 1685 3507 1686 3559
rect 1632 3506 1686 3507
rect 1632 3071 1686 3072
rect 1632 3019 1633 3071
rect 1685 3019 1686 3071
rect 1632 3018 1686 3019
rect 3802 3051 3838 3052
rect 3802 3017 3803 3051
rect 3837 3017 3838 3051
rect 3802 3016 3838 3017
rect 3894 3051 3930 3052
rect 3894 3017 3895 3051
rect 3929 3017 3930 3051
rect 3894 3016 3930 3017
rect 40 2993 76 2994
rect 40 2959 41 2993
rect 75 2959 76 2993
rect 40 2958 76 2959
rect 132 2993 168 2994
rect 132 2959 133 2993
rect 167 2959 168 2993
rect 132 2958 168 2959
rect 1632 2971 1686 2972
rect 1632 2919 1633 2971
rect 1685 2919 1686 2971
rect 3802 2959 3838 2960
rect 3802 2925 3803 2959
rect 3837 2925 3838 2959
rect 3802 2924 3838 2925
rect 3894 2959 3930 2960
rect 3894 2925 3895 2959
rect 3929 2925 3930 2959
rect 3894 2924 3930 2925
rect 1632 2918 1686 2919
rect 1632 2623 1686 2624
rect 1632 2571 1633 2623
rect 1685 2571 1686 2623
rect 1632 2570 1686 2571
rect 3802 2591 3838 2592
rect 3802 2564 3803 2591
rect 16 2533 184 2564
rect 16 2530 41 2533
rect 40 2499 41 2530
rect 75 2530 133 2533
rect 75 2499 76 2530
rect 40 2498 76 2499
rect 132 2499 133 2530
rect 167 2530 184 2533
rect 3774 2557 3803 2564
rect 3837 2564 3838 2591
rect 3894 2591 3930 2592
rect 3894 2564 3895 2591
rect 3837 2557 3895 2564
rect 3929 2564 3930 2591
rect 3929 2557 3946 2564
rect 167 2499 168 2530
rect 132 2498 168 2499
rect 1632 2523 1686 2524
rect 1632 2471 1633 2523
rect 1685 2471 1686 2523
rect 3774 2499 3946 2557
rect 3774 2486 3803 2499
rect 1632 2470 1686 2471
rect 3802 2465 3803 2486
rect 3837 2486 3895 2499
rect 3837 2465 3838 2486
rect 3802 2464 3838 2465
rect 3894 2465 3895 2486
rect 3929 2486 3946 2499
rect 3929 2465 3930 2486
rect 3894 2464 3930 2465
rect 1632 2179 1686 2180
rect 1632 2127 1633 2179
rect 1685 2127 1686 2179
rect 1632 2126 1686 2127
rect 3774 2131 3946 2164
rect 16 2086 184 2120
rect 3774 2097 3803 2131
rect 3837 2097 3895 2131
rect 3929 2097 3946 2131
rect 3774 2086 3946 2097
rect 1632 2079 1686 2080
rect 1632 2027 1633 2079
rect 1685 2027 1686 2079
rect 1632 2026 1686 2027
rect 1632 1415 1686 1416
rect 1632 1363 1633 1415
rect 1685 1363 1686 1415
rect 1632 1362 1686 1363
rect 3802 1395 3838 1396
rect 3802 1361 3803 1395
rect 3837 1361 3838 1395
rect 3802 1360 3838 1361
rect 3894 1395 3930 1396
rect 3894 1361 3895 1395
rect 3929 1361 3930 1395
rect 3894 1360 3930 1361
rect 1632 1315 1686 1316
rect 1632 1263 1633 1315
rect 1685 1263 1686 1315
rect 3802 1303 3838 1304
rect 3802 1269 3803 1303
rect 3837 1269 3838 1303
rect 3802 1268 3838 1269
rect 1632 1262 1686 1263
rect 1634 59 1688 60
rect 1634 7 1635 59
rect 1687 7 1688 59
rect 1634 6 1688 7
<< via1 >>
rect 1633 5027 1685 5079
rect 1633 4235 1685 4287
rect 1633 4115 1685 4167
rect 1633 3627 1685 3679
rect 1633 3507 1685 3559
rect 1633 3019 1685 3071
rect 1633 2919 1685 2971
rect 1633 2571 1685 2623
rect 1633 2471 1685 2523
rect 1633 2127 1685 2179
rect 1633 2027 1685 2079
rect 1633 1363 1685 1415
rect 1633 1263 1685 1315
rect 1635 7 1687 59
<< metal2 >>
rect 1626 5079 1692 5086
rect 1626 5027 1633 5079
rect 1685 5070 1692 5079
rect 1685 5036 1756 5070
rect 1685 5027 1692 5036
rect 1626 5020 1692 5027
rect 1626 4287 1692 4294
rect 1626 4235 1633 4287
rect 1685 4235 1692 4287
rect 1626 4228 1692 4235
rect 1626 4167 1692 4174
rect 1626 4115 1633 4167
rect 1685 4158 1692 4167
rect 1722 4158 1756 5036
rect 1685 4124 1756 4158
rect 1685 4115 1692 4124
rect 1626 4108 1692 4115
rect 1626 3679 1692 3686
rect 1626 3627 1633 3679
rect 1685 3627 1692 3679
rect 1626 3620 1692 3627
rect 1626 3559 1692 3566
rect 1626 3507 1633 3559
rect 1685 3550 1692 3559
rect 1722 3550 1756 4124
rect 1685 3516 1756 3550
rect 1685 3507 1692 3516
rect 1626 3500 1692 3507
rect 1626 3071 1692 3078
rect 1626 3019 1633 3071
rect 1685 3019 1692 3071
rect 1626 3012 1692 3019
rect 1626 2971 1692 2978
rect 1626 2919 1633 2971
rect 1685 2962 1692 2971
rect 1722 2962 1756 3516
rect 1685 2928 1756 2962
rect 1685 2919 1692 2928
rect 1626 2912 1692 2919
rect 1626 2623 1692 2630
rect 1626 2571 1633 2623
rect 1685 2571 1692 2623
rect 1626 2564 1692 2571
rect 1626 2523 1692 2530
rect 1626 2471 1633 2523
rect 1685 2514 1692 2523
rect 1722 2514 1756 2928
rect 1685 2480 1756 2514
rect 1685 2471 1692 2480
rect 1626 2464 1692 2471
rect 1626 2179 1692 2186
rect 1626 2127 1633 2179
rect 1685 2127 1692 2179
rect 1626 2120 1692 2127
rect 1626 2079 1692 2086
rect 1626 2027 1633 2079
rect 1685 2070 1692 2079
rect 1722 2070 1756 2480
rect 1685 2036 1756 2070
rect 1685 2027 1692 2036
rect 1626 2020 1692 2027
rect 1626 1415 1692 1422
rect 1626 1363 1633 1415
rect 1685 1363 1692 1415
rect 1626 1356 1692 1363
rect 1626 1315 1692 1322
rect 1626 1263 1633 1315
rect 1685 1306 1692 1315
rect 1722 1306 1756 2036
rect 1685 1272 1756 1306
rect 1685 1263 1692 1272
rect 1626 1256 1692 1263
rect 1628 59 1694 66
rect 1628 7 1635 59
rect 1687 7 1694 59
rect 1628 0 1694 7
use inverter_p0o47_n40  inverter_p0o47_n40_0
timestamp 1756008383
transform 0 1 166 -1 0 5086
box -62 -192 920 3830
use inverter_p2_n18  inverter_p2_n18_0
timestamp 1756008383
transform 0 1 600 -1 0 4174
box -36 -626 616 3396
use inverter_p7_n10  inverter_p7_n10_0
timestamp 1756008383
transform 0 1 1000 -1 0 3566
box -142 -1026 590 3128
use inverter_p15_n5  inverter_p15_n5_0
timestamp 1756008383
transform 0 1 1000 -1 0 2898
box -108 -1026 360 2996
use inverter_p16_n1o5  inverter_p16_n1o5_0
timestamp 1756008383
transform 0 1 1262 -1 0 2442
box -114 -1288 474 2734
use inverter_p40_n1  inverter_p40_n1_0
timestamp 1756008383
transform 0 1 1350 -1 0 1838
box -274 -1376 634 2646
use inverter_p90_n0o47  inverter_p90_n0o47_0
timestamp 1756008383
transform 0 1 1456 -1 0 730
box -664 -1482 756 2540
<< end >>
