magic
tech sky130A
magscale 1 2
timestamp 1752540706
<< nwell >>
rect -36 544 182 674
<< psubdiff >>
rect 2 -52 148 -32
rect 2 -86 28 -52
rect 124 -86 148 -52
rect 2 -106 148 -86
<< nsubdiff >>
rect 0 604 146 620
rect 0 570 40 604
rect 106 570 146 604
rect 0 546 146 570
<< psubdiffcont >>
rect 28 -86 124 -52
<< nsubdiffcont >>
rect 40 570 106 604
<< poly >>
rect 58 226 88 276
rect -8 210 88 226
rect -8 176 8 210
rect 42 176 88 210
rect -8 162 88 176
rect 58 136 88 162
<< polycont >>
rect 8 176 42 210
<< locali >>
rect 6 604 140 614
rect 6 570 40 604
rect 106 570 140 604
rect 6 552 140 570
rect 12 486 46 552
rect 100 226 134 298
rect -36 210 58 226
rect -36 176 8 210
rect 42 176 58 210
rect -36 162 58 176
rect 100 164 182 226
rect 100 114 134 164
rect 12 -40 46 22
rect 10 -52 140 -40
rect 10 -86 28 -52
rect 124 -86 140 -52
rect 10 -98 140 -86
<< viali >>
rect 40 570 106 604
rect 28 -86 124 -52
<< metal1 >>
rect -36 604 182 614
rect -36 570 40 604
rect 106 570 182 604
rect -36 552 182 570
rect 12 470 46 552
rect 10 -40 46 38
rect -34 -52 182 -40
rect -34 -86 28 -52
rect 124 -86 182 -52
rect -34 -98 182 -86
use sky130_fd_pr__nfet_01v8_HEP5MT  sky130_fd_pr__nfet_01v8_HEP5MT_0
timestamp 1752539806
transform 1 0 73 0 1 68
box -73 -68 73 68
use sky130_fd_pr__pfet_01v8_35B5V5  sky130_fd_pr__pfet_01v8_35B5V5_0
timestamp 1752539806
transform 1 0 73 0 1 392
box -109 -152 109 152
<< labels >>
rlabel locali -26 202 -26 202 7 Vin
port 1 w
rlabel locali 178 198 178 198 3 Vout
port 2 e
rlabel metal1 6 584 6 584 7 VDD
port 3 w
rlabel metal1 10 -68 10 -68 7 GND
port 4 w
<< end >>
