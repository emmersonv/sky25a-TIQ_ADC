magic
tech sky130A
timestamp 1755919380
<< nwell >>
rect 861 2508 878 2518
rect 1880 2105 1980 2115
rect 1117 1801 1998 2105
rect 1880 1783 1980 1801
rect 1901 1508 1919 1526
rect 1947 1508 1965 1526
rect 861 1282 878 1464
rect 1880 1449 1980 1506
rect 1880 1282 1980 1323
rect 828 1243 1998 1282
rect 1880 1225 1980 1243
rect 1880 1082 1980 1100
rect 822 1017 1998 1082
rect 1880 999 1980 1017
rect 1880 704 1980 722
rect 822 635 1998 704
rect 1880 617 1980 635
<< psubdiff >>
rect 0 2095 100 2096
rect 0 2087 20 2095
rect 38 2087 66 2095
rect 84 2087 100 2095
rect 0 1783 100 1792
rect 0 1497 100 1506
rect 0 1490 20 1497
rect 38 1490 66 1497
rect 84 1490 100 1497
rect 0 1267 100 1282
rect 0 1265 20 1267
rect 38 1265 66 1267
rect 84 1265 100 1267
rect 0 1043 100 1060
<< nsubdiff >>
rect 1880 2087 1980 2115
rect 1880 1802 1980 1810
rect 1880 1784 1901 1802
rect 1919 1784 1947 1802
rect 1965 1784 1980 1802
rect 1880 1783 1980 1784
rect 1880 1480 1980 1506
rect 1880 1462 1901 1480
rect 1919 1462 1947 1480
rect 1965 1462 1980 1480
rect 1880 1449 1980 1462
rect 1880 1296 1980 1323
rect 1880 1278 1901 1296
rect 1919 1278 1947 1296
rect 1965 1278 1980 1296
rect 1880 1250 1980 1278
rect 1880 1232 1901 1250
rect 1919 1232 1947 1250
rect 1965 1232 1980 1250
rect 1880 1225 1980 1232
rect 1880 1094 1901 1100
rect 1919 1094 1947 1100
rect 1965 1094 1980 1100
rect 1880 1066 1980 1094
rect 1880 1048 1901 1066
rect 1919 1048 1947 1066
rect 1965 1048 1980 1066
rect 1880 1020 1980 1048
rect 1880 1002 1901 1020
rect 1919 1002 1947 1020
rect 1965 1002 1980 1020
rect 1880 999 1980 1002
rect 1880 698 1980 722
rect 1880 680 1901 698
rect 1919 680 1947 698
rect 1965 680 1980 698
rect 1880 652 1980 680
rect 1880 634 1901 652
rect 1919 634 1947 652
rect 1965 634 1980 652
rect 1880 617 1980 634
<< psubdiffcont >>
rect 20 2077 38 2095
rect 66 2077 84 2095
rect 20 1479 38 1497
rect 66 1479 84 1497
rect 20 1249 38 1267
rect 66 1249 84 1267
<< nsubdiffcont >>
rect 1901 1784 1919 1802
rect 1947 1784 1965 1802
rect 1901 1508 1919 1526
rect 1947 1508 1965 1526
rect 1901 1462 1919 1480
rect 1947 1462 1965 1480
rect 1901 1324 1919 1342
rect 1947 1324 1965 1342
rect 1901 1278 1919 1296
rect 1947 1278 1965 1296
rect 1901 1232 1919 1250
rect 1947 1232 1965 1250
rect 1901 1094 1919 1112
rect 1947 1094 1965 1112
rect 1901 1048 1919 1066
rect 1947 1048 1965 1066
rect 1901 1002 1919 1020
rect 1947 1002 1965 1020
rect 1901 680 1919 698
rect 1947 680 1965 698
rect 1901 634 1919 652
rect 1947 634 1965 652
<< locali >>
rect 8 2095 92 2096
rect 8 2087 20 2095
rect 38 2087 66 2095
rect 84 2087 92 2095
rect 8 1267 92 1282
rect 8 1265 20 1267
rect 38 1265 66 1267
rect 84 1265 92 1267
rect 1887 1278 1901 1282
rect 1919 1278 1947 1282
rect 1965 1278 1973 1282
rect 1887 1250 1973 1278
rect 1887 1243 1901 1250
rect 1919 1243 1947 1250
rect 1965 1243 1973 1250
rect 1887 1066 1973 1082
rect 8 1043 92 1060
rect 1887 1048 1901 1066
rect 1919 1048 1947 1066
rect 1965 1048 1973 1066
rect 1887 1043 1973 1048
<< viali >>
rect 20 2077 38 2095
rect 66 2077 84 2095
rect 1901 1784 1919 1802
rect 1947 1784 1965 1802
rect 1901 1508 1919 1526
rect 1947 1508 1965 1526
rect 20 1479 38 1497
rect 66 1479 84 1497
rect 1901 1462 1919 1480
rect 1947 1462 1965 1480
rect 20 1249 38 1267
rect 66 1249 84 1267
rect 1901 1278 1919 1296
rect 1947 1278 1965 1296
rect 1901 1232 1919 1250
rect 1947 1232 1965 1250
rect 1901 1048 1919 1066
rect 1947 1048 1965 1066
rect 1901 680 1919 698
rect 1947 680 1965 698
rect 1901 634 1919 652
<< metal1 >>
rect 8 2095 92 2096
rect 8 2087 20 2095
rect 38 2087 66 2095
rect 84 2087 92 2095
rect 8 1267 92 1282
rect 8 1265 20 1267
rect 38 1265 66 1267
rect 84 1265 92 1267
rect 1887 1278 1901 1282
rect 1919 1278 1947 1282
rect 1965 1278 1973 1282
rect 1887 1250 1973 1278
rect 1887 1243 1901 1250
rect 1919 1243 1947 1250
rect 1965 1243 1973 1250
rect 1887 1066 1973 1082
rect 8 1043 92 1060
rect 1887 1048 1901 1066
rect 1919 1048 1947 1066
rect 1965 1048 1973 1066
rect 1887 1043 1973 1048
<< via1 >>
rect 816 2513 843 2540
rect 816 2117 843 2144
rect 816 2057 843 2084
rect 816 1813 843 1840
rect 816 1753 843 1780
rect 816 1509 843 1536
rect 816 1459 843 1486
rect 816 1285 843 1312
rect 816 1235 843 1262
rect 816 1063 843 1090
rect 816 1013 843 1040
rect 816 681 843 708
rect 816 631 843 658
rect 817 3 844 30
<< metal2 >>
rect 813 2540 846 2543
rect 813 2513 816 2540
rect 843 2535 846 2540
rect 843 2518 878 2535
rect 843 2513 846 2518
rect 813 2510 846 2513
rect 813 2144 846 2147
rect 813 2117 816 2144
rect 843 2117 846 2144
rect 813 2114 846 2117
rect 813 2084 846 2087
rect 813 2057 816 2084
rect 843 2079 846 2084
rect 861 2079 878 2518
rect 843 2062 878 2079
rect 843 2057 846 2062
rect 813 2054 846 2057
rect 813 1840 846 1843
rect 813 1813 816 1840
rect 843 1813 846 1840
rect 813 1810 846 1813
rect 813 1780 846 1783
rect 813 1753 816 1780
rect 843 1775 846 1780
rect 861 1775 878 2062
rect 843 1758 878 1775
rect 843 1753 846 1758
rect 813 1750 846 1753
rect 813 1536 846 1539
rect 813 1509 816 1536
rect 843 1509 846 1536
rect 813 1506 846 1509
rect 813 1486 846 1489
rect 813 1459 816 1486
rect 843 1481 846 1486
rect 861 1481 878 1758
rect 843 1464 878 1481
rect 843 1459 846 1464
rect 813 1456 846 1459
rect 813 1312 846 1315
rect 813 1285 816 1312
rect 843 1285 846 1312
rect 813 1282 846 1285
rect 813 1262 846 1265
rect 813 1235 816 1262
rect 843 1257 846 1262
rect 861 1257 878 1464
rect 843 1240 878 1257
rect 843 1235 846 1240
rect 813 1232 846 1235
rect 813 1090 846 1093
rect 813 1063 816 1090
rect 843 1063 846 1090
rect 813 1060 846 1063
rect 813 1040 846 1043
rect 813 1013 816 1040
rect 843 1035 846 1040
rect 861 1035 878 1240
rect 843 1018 878 1035
rect 843 1013 846 1018
rect 813 1010 846 1013
rect 813 708 846 711
rect 813 681 816 708
rect 843 681 846 708
rect 813 678 846 681
rect 813 658 846 661
rect 813 631 816 658
rect 843 653 846 658
rect 861 653 878 1018
rect 843 636 878 653
rect 843 631 846 636
rect 813 628 846 631
rect 814 30 847 33
rect 814 3 817 30
rect 844 3 847 30
rect 814 0 847 3
use inverter_p0o47_n40  inverter_p0o47_n40_0
timestamp 1755919380
transform 0 1 83 -1 0 2543
box -18 -83 447 1915
use inverter_p2_n18  inverter_p2_n18_0
timestamp 1755919380
transform 0 1 300 -1 0 2087
box -18 -300 367 1698
use inverter_p7_n10  inverter_p7_n10_0
timestamp 1755919380
transform 0 1 500 -1 0 1783
box -18 -500 295 1498
use inverter_p15_n5  inverter_p15_n5_0
timestamp 1755919380
transform 0 1 500 -1 0 1449
box -41 -500 167 1498
use inverter_p16_n1o5  inverter_p16_n1o5_0
timestamp 1755919380
transform 0 1 631 -1 0 1221
box -44 -631 237 1367
use inverter_p40_n1  inverter_p40_n1_0
timestamp 1755919380
transform 0 1 675 -1 0 919
box -124 -675 317 1323
use inverter_p90_n0o47  inverter_p90_n0o47_0
timestamp 1755919380
transform 0 1 728 -1 0 365
box -319 -728 365 1270
<< end >>
