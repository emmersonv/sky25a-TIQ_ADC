magic
tech sky130A
magscale 1 2
timestamp 1756008383
<< pwell >>
rect -99 -68 99 68
<< nmos >>
rect -15 -42 15 42
<< ndiff >>
rect -73 17 -15 42
rect -73 -17 -61 17
rect -27 -17 -15 17
rect -73 -42 -15 -17
rect 15 17 73 42
rect 15 -17 27 17
rect 61 -17 73 17
rect 15 -42 73 -17
<< ndiffc >>
rect -61 -17 -27 17
rect 27 -17 61 17
<< poly >>
rect -15 42 15 68
rect -15 -68 15 -42
<< locali >>
rect -61 17 -27 46
rect -61 -46 -27 -17
rect 27 17 61 46
rect 27 -46 61 -17
<< viali >>
rect -61 -17 -27 17
rect 27 -17 61 17
<< metal1 >>
rect -67 17 -21 42
rect -67 -17 -61 17
rect -27 -17 -21 17
rect -67 -42 -21 -17
rect 21 17 67 42
rect 21 -17 27 17
rect 61 -17 67 17
rect 21 -42 67 -17
<< end >>
