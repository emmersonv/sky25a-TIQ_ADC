magic
tech sky130A
magscale 1 2
timestamp 1756008383
<< pwell >>
rect -99 -176 99 176
<< nmos >>
rect -15 -150 15 150
<< ndiff >>
rect -73 119 -15 150
rect -73 85 -61 119
rect -27 85 -15 119
rect -73 51 -15 85
rect -73 17 -61 51
rect -27 17 -15 51
rect -73 -17 -15 17
rect -73 -51 -61 -17
rect -27 -51 -15 -17
rect -73 -85 -15 -51
rect -73 -119 -61 -85
rect -27 -119 -15 -85
rect -73 -150 -15 -119
rect 15 119 73 150
rect 15 85 27 119
rect 61 85 73 119
rect 15 51 73 85
rect 15 17 27 51
rect 61 17 73 51
rect 15 -17 73 17
rect 15 -51 27 -17
rect 61 -51 73 -17
rect 15 -85 73 -51
rect 15 -119 27 -85
rect 61 -119 73 -85
rect 15 -150 73 -119
<< ndiffc >>
rect -61 85 -27 119
rect -61 17 -27 51
rect -61 -51 -27 -17
rect -61 -119 -27 -85
rect 27 85 61 119
rect 27 17 61 51
rect 27 -51 61 -17
rect 27 -119 61 -85
<< poly >>
rect -15 150 15 176
rect -15 -176 15 -150
<< locali >>
rect -61 125 -27 154
rect -61 53 -27 85
rect -61 -17 -27 17
rect -61 -85 -27 -53
rect -61 -154 -27 -125
rect 27 125 61 154
rect 27 53 61 85
rect 27 -17 61 17
rect 27 -85 61 -53
rect 27 -154 61 -125
<< viali >>
rect -61 119 -27 125
rect -61 91 -27 119
rect -61 51 -27 53
rect -61 19 -27 51
rect -61 -51 -27 -19
rect -61 -53 -27 -51
rect -61 -119 -27 -91
rect -61 -125 -27 -119
rect 27 119 61 125
rect 27 91 61 119
rect 27 51 61 53
rect 27 19 61 51
rect 27 -51 61 -19
rect 27 -53 61 -51
rect 27 -119 61 -91
rect 27 -125 61 -119
<< metal1 >>
rect -67 125 -21 150
rect -67 91 -61 125
rect -27 91 -21 125
rect -67 53 -21 91
rect -67 19 -61 53
rect -27 19 -21 53
rect -67 -19 -21 19
rect -67 -53 -61 -19
rect -27 -53 -21 -19
rect -67 -91 -21 -53
rect -67 -125 -61 -91
rect -27 -125 -21 -91
rect -67 -150 -21 -125
rect 21 125 67 150
rect 21 91 27 125
rect 61 91 67 125
rect 21 53 67 91
rect 21 19 27 53
rect 61 19 67 53
rect 21 -19 67 19
rect 21 -53 27 -19
rect 61 -53 67 -19
rect 21 -91 67 -53
rect 21 -125 27 -91
rect 61 -125 67 -91
rect 21 -150 67 -125
<< end >>
