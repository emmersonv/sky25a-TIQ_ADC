magic
tech sky130A
magscale 1 2
timestamp 1756008383
<< pwell >>
rect -151 -276 151 276
<< nmos >>
rect -63 -250 -33 250
rect 33 -250 63 250
<< ndiff >>
rect -125 221 -63 250
rect -125 187 -113 221
rect -79 187 -63 221
rect -125 153 -63 187
rect -125 119 -113 153
rect -79 119 -63 153
rect -125 85 -63 119
rect -125 51 -113 85
rect -79 51 -63 85
rect -125 17 -63 51
rect -125 -17 -113 17
rect -79 -17 -63 17
rect -125 -51 -63 -17
rect -125 -85 -113 -51
rect -79 -85 -63 -51
rect -125 -119 -63 -85
rect -125 -153 -113 -119
rect -79 -153 -63 -119
rect -125 -187 -63 -153
rect -125 -221 -113 -187
rect -79 -221 -63 -187
rect -125 -250 -63 -221
rect -33 221 33 250
rect -33 187 -17 221
rect 17 187 33 221
rect -33 153 33 187
rect -33 119 -17 153
rect 17 119 33 153
rect -33 85 33 119
rect -33 51 -17 85
rect 17 51 33 85
rect -33 17 33 51
rect -33 -17 -17 17
rect 17 -17 33 17
rect -33 -51 33 -17
rect -33 -85 -17 -51
rect 17 -85 33 -51
rect -33 -119 33 -85
rect -33 -153 -17 -119
rect 17 -153 33 -119
rect -33 -187 33 -153
rect -33 -221 -17 -187
rect 17 -221 33 -187
rect -33 -250 33 -221
rect 63 221 125 250
rect 63 187 79 221
rect 113 187 125 221
rect 63 153 125 187
rect 63 119 79 153
rect 113 119 125 153
rect 63 85 125 119
rect 63 51 79 85
rect 113 51 125 85
rect 63 17 125 51
rect 63 -17 79 17
rect 113 -17 125 17
rect 63 -51 125 -17
rect 63 -85 79 -51
rect 113 -85 125 -51
rect 63 -119 125 -85
rect 63 -153 79 -119
rect 113 -153 125 -119
rect 63 -187 125 -153
rect 63 -221 79 -187
rect 113 -221 125 -187
rect 63 -250 125 -221
<< ndiffc >>
rect -113 187 -79 221
rect -113 119 -79 153
rect -113 51 -79 85
rect -113 -17 -79 17
rect -113 -85 -79 -51
rect -113 -153 -79 -119
rect -113 -221 -79 -187
rect -17 187 17 221
rect -17 119 17 153
rect -17 51 17 85
rect -17 -17 17 17
rect -17 -85 17 -51
rect -17 -153 17 -119
rect -17 -221 17 -187
rect 79 187 113 221
rect 79 119 113 153
rect 79 51 113 85
rect 79 -17 113 17
rect 79 -85 113 -51
rect 79 -153 113 -119
rect 79 -221 113 -187
<< poly >>
rect -63 276 63 306
rect -63 250 -33 276
rect 33 250 63 276
rect -63 -276 -33 -250
rect 33 -276 63 -250
<< locali >>
rect -113 233 -79 254
rect -113 161 -79 187
rect -113 89 -79 119
rect -113 17 -79 51
rect -113 -51 -79 -17
rect -113 -119 -79 -89
rect -113 -187 -79 -161
rect -113 -254 -79 -233
rect -17 233 17 254
rect -17 161 17 187
rect -17 89 17 119
rect -17 17 17 51
rect -17 -51 17 -17
rect -17 -119 17 -89
rect -17 -187 17 -161
rect -17 -254 17 -233
rect 79 233 113 254
rect 79 161 113 187
rect 79 89 113 119
rect 79 17 113 51
rect 79 -51 113 -17
rect 79 -119 113 -89
rect 79 -187 113 -161
rect 79 -254 113 -233
<< viali >>
rect -113 221 -79 233
rect -113 199 -79 221
rect -113 153 -79 161
rect -113 127 -79 153
rect -113 85 -79 89
rect -113 55 -79 85
rect -113 -17 -79 17
rect -113 -85 -79 -55
rect -113 -89 -79 -85
rect -113 -153 -79 -127
rect -113 -161 -79 -153
rect -113 -221 -79 -199
rect -113 -233 -79 -221
rect -17 221 17 233
rect -17 199 17 221
rect -17 153 17 161
rect -17 127 17 153
rect -17 85 17 89
rect -17 55 17 85
rect -17 -17 17 17
rect -17 -85 17 -55
rect -17 -89 17 -85
rect -17 -153 17 -127
rect -17 -161 17 -153
rect -17 -221 17 -199
rect -17 -233 17 -221
rect 79 221 113 233
rect 79 199 113 221
rect 79 153 113 161
rect 79 127 113 153
rect 79 85 113 89
rect 79 55 113 85
rect 79 -17 113 17
rect 79 -85 113 -55
rect 79 -89 113 -85
rect 79 -153 113 -127
rect 79 -161 113 -153
rect 79 -221 113 -199
rect 79 -233 113 -221
<< metal1 >>
rect -119 233 -73 250
rect -119 199 -113 233
rect -79 199 -73 233
rect -119 161 -73 199
rect -119 127 -113 161
rect -79 127 -73 161
rect -119 89 -73 127
rect -119 55 -113 89
rect -79 55 -73 89
rect -119 17 -73 55
rect -119 -17 -113 17
rect -79 -17 -73 17
rect -119 -55 -73 -17
rect -119 -89 -113 -55
rect -79 -89 -73 -55
rect -119 -127 -73 -89
rect -119 -161 -113 -127
rect -79 -161 -73 -127
rect -119 -199 -73 -161
rect -119 -233 -113 -199
rect -79 -233 -73 -199
rect -119 -250 -73 -233
rect -23 233 23 250
rect -23 199 -17 233
rect 17 199 23 233
rect -23 161 23 199
rect -23 127 -17 161
rect 17 127 23 161
rect -23 89 23 127
rect -23 55 -17 89
rect 17 55 23 89
rect -23 17 23 55
rect -23 -17 -17 17
rect 17 -17 23 17
rect -23 -55 23 -17
rect -23 -89 -17 -55
rect 17 -89 23 -55
rect -23 -127 23 -89
rect -23 -161 -17 -127
rect 17 -161 23 -127
rect -23 -199 23 -161
rect -23 -233 -17 -199
rect 17 -233 23 -199
rect -23 -250 23 -233
rect 73 233 119 250
rect 73 199 79 233
rect 113 199 119 233
rect 73 161 119 199
rect 73 127 79 161
rect 113 127 119 161
rect 73 89 119 127
rect 73 55 79 89
rect 113 55 119 89
rect 73 17 119 55
rect 73 -17 79 17
rect 113 -17 119 17
rect 73 -55 119 -17
rect 73 -89 79 -55
rect 113 -89 119 -55
rect 73 -127 119 -89
rect 73 -161 79 -127
rect 113 -161 119 -127
rect 73 -199 119 -161
rect 73 -233 79 -199
rect 113 -233 119 -199
rect 73 -250 119 -233
<< end >>
