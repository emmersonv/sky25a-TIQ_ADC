magic
tech sky130A
magscale 1 2
timestamp 1754101402
<< error_p >>
rect -125 -250 -63 250
rect -33 -250 33 250
rect 63 -250 125 250
<< nmos >>
rect -63 -250 -33 250
rect 33 -250 63 250
<< ndiff >>
rect -125 238 -63 250
rect -125 -238 -113 238
rect -79 -238 -63 238
rect -125 -250 -63 -238
rect -33 238 33 250
rect -33 -238 -17 238
rect 17 -238 33 238
rect -33 -250 33 -238
rect 63 238 125 250
rect 63 -238 79 238
rect 113 -238 125 238
rect 63 -250 125 -238
<< ndiffc >>
rect -113 -238 -79 238
rect -17 -238 17 238
rect 79 -238 113 238
<< poly >>
rect -63 276 63 306
rect -63 250 -33 276
rect 33 250 63 276
rect -63 -276 -33 -250
rect 33 -276 63 -250
<< locali >>
rect -113 238 -79 254
rect -113 -254 -79 -238
rect -17 238 17 254
rect -17 -254 17 -238
rect 79 238 113 254
rect 79 -254 113 -238
<< viali >>
rect -113 -238 -79 238
rect -17 -238 17 238
rect 79 -238 113 238
<< metal1 >>
rect -119 238 -73 250
rect -119 -238 -113 238
rect -79 -238 -73 238
rect -119 -250 -73 -238
rect -23 238 23 250
rect -23 -238 -17 238
rect 17 -238 23 238
rect -23 -250 23 -238
rect 73 238 119 250
rect 73 -238 79 238
rect 113 -238 119 238
rect 73 -250 119 -238
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 2.5 l 0.150 m 1 nf 2 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 class mosfet compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
