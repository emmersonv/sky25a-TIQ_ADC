* NGSPICE file created from inverter_p1_n15.ext - technology: sky130A

.subckt sky130_fd_pr__pfet_01v8_TH65V5 a_n73_n100# w_n109_n162# a_15_n100# a_n15_n126#
X0 a_15_n100# a_n15_n126# a_n73_n100# w_n109_n162# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
.ends

.subckt sky130_fd_pr__nfet_01v8_3LPVTD a_63_n750# a_n63_n776# a_n33_n750# a_n125_n750#
+ VSUBS
X0 a_63_n750# a_n63_n776# a_n33_n750# VSUBS sky130_fd_pr__nfet_01v8 ad=2.325 pd=15.62 as=1.2375 ps=7.83 w=7.5 l=0.15
X1 a_n33_n750# a_n63_n776# a_n125_n750# VSUBS sky130_fd_pr__nfet_01v8 ad=1.2375 pd=7.83 as=2.325 ps=15.62 w=7.5 l=0.15
.ends

.subckt inverter_p1_n15 VDPWR Vout Vin VGND
Xsky130_fd_pr__pfet_01v8_TH65V5_0 VDPWR VDPWR Vout Vin sky130_fd_pr__pfet_01v8_TH65V5
Xsky130_fd_pr__nfet_01v8_3LPVTD_0 VGND Vin Vout VGND VGND sky130_fd_pr__nfet_01v8_3LPVTD
.ends

