magic
tech sky130A
magscale 1 2
timestamp 1754112194
<< nwell >>
rect -80 656 334 2996
<< psubdiff >>
rect -82 -832 334 -800
rect -82 -868 -4 -832
rect 32 -868 88 -832
rect 124 -868 180 -832
rect 216 -868 272 -832
rect 308 -868 334 -832
rect -82 -924 334 -868
rect -82 -960 -4 -924
rect 32 -960 88 -924
rect 124 -960 180 -924
rect 216 -960 272 -924
rect 308 -960 334 -924
rect -82 -1000 334 -960
<< nsubdiff >>
rect 0 2930 252 2960
rect 0 2894 30 2930
rect 66 2894 122 2930
rect 158 2894 252 2930
rect 0 2838 252 2894
rect 0 2802 30 2838
rect 66 2802 122 2838
rect 158 2802 252 2838
rect 0 2760 252 2802
<< psubdiffcont >>
rect -4 -868 32 -832
rect 88 -868 124 -832
rect 180 -868 216 -832
rect 272 -868 308 -832
rect -4 -960 32 -924
rect 88 -960 124 -924
rect 180 -960 216 -924
rect 272 -960 308 -924
<< nsubdiffcont >>
rect 30 2894 66 2930
rect 122 2894 158 2930
rect 30 2802 66 2838
rect 122 2802 158 2838
<< poly >>
rect -80 676 -14 692
rect -80 642 -64 676
rect -30 656 -14 676
rect 62 656 188 662
rect -30 644 188 656
rect -30 642 62 644
rect -80 626 62 642
<< polycont >>
rect -64 642 -30 676
<< locali >>
rect -80 2930 334 2946
rect -80 2894 -62 2930
rect -26 2894 30 2930
rect 66 2894 122 2930
rect 158 2894 214 2930
rect 250 2894 334 2930
rect -80 2838 334 2894
rect -80 2802 -62 2838
rect -26 2802 30 2838
rect 66 2802 122 2838
rect 158 2802 214 2838
rect 250 2802 334 2838
rect -80 2774 334 2802
rect 12 2222 46 2774
rect 204 2222 238 2774
rect -80 676 -14 692
rect -80 642 -64 676
rect -30 642 -14 676
rect -80 626 -14 642
rect 108 666 142 714
rect 268 676 334 692
rect 268 666 284 676
rect 108 642 284 666
rect 318 642 334 676
rect 108 626 334 642
rect 108 592 142 626
rect 12 -816 46 84
rect 204 -816 238 84
rect -80 -832 334 -816
rect -80 -868 -4 -832
rect 32 -868 88 -832
rect 124 -868 180 -832
rect 216 -868 272 -832
rect 308 -868 334 -832
rect -80 -924 334 -868
rect -80 -960 -4 -924
rect 32 -960 88 -924
rect 124 -960 180 -924
rect 216 -960 272 -924
rect 308 -960 334 -924
rect -80 -984 334 -960
<< viali >>
rect -62 2894 -26 2930
rect 30 2894 66 2930
rect 122 2894 158 2930
rect 214 2894 250 2930
rect -62 2802 -26 2838
rect 30 2802 66 2838
rect 122 2802 158 2838
rect 214 2802 250 2838
rect -64 642 -30 676
rect 284 642 318 676
rect -4 -868 32 -832
rect 88 -868 124 -832
rect 180 -868 216 -832
rect 272 -868 308 -832
rect -4 -960 32 -924
rect 88 -960 124 -924
rect 180 -960 216 -924
rect 272 -960 308 -924
<< metal1 >>
rect -80 2930 334 2946
rect -80 2894 -62 2930
rect -26 2894 30 2930
rect 66 2894 122 2930
rect 158 2894 214 2930
rect 250 2894 334 2930
rect -80 2838 334 2894
rect -80 2802 -62 2838
rect -26 2802 30 2838
rect 66 2802 122 2838
rect 158 2802 214 2838
rect 250 2802 334 2838
rect -80 2774 334 2802
rect -80 676 -14 692
rect -80 642 -64 676
rect -30 642 -14 676
rect -80 626 -14 642
rect 268 676 334 692
rect 268 642 284 676
rect 318 642 334 676
rect 268 626 334 642
rect -80 -832 334 -816
rect -80 -868 -4 -832
rect 32 -868 88 -832
rect 124 -868 180 -832
rect 216 -868 272 -832
rect 308 -868 334 -832
rect -80 -924 334 -868
rect -80 -960 -4 -924
rect 32 -960 88 -924
rect 124 -960 180 -924
rect 216 -960 272 -924
rect 308 -960 334 -924
rect -80 -984 334 -960
use sky130_fd_pr__nfet_01v8_V2VUT3  sky130_fd_pr__nfet_01v8_V2VUT3_0
timestamp 1754101402
transform 1 0 125 0 1 338
box -125 -276 125 306
use sky130_fd_pr__pfet_01v8_7QKTNL  sky130_fd_pr__pfet_01v8_7QKTNL_0
timestamp 1753684791
transform 1 0 125 0 1 1468
box -161 -812 161 812
<< end >>
