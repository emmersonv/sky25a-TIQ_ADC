magic
tech sky130A
magscale 1 2
timestamp 1755919380
<< viali >>
rect 6285 6205 6319 6239
rect 6561 6205 6595 6239
rect 6101 6069 6135 6103
rect 6377 6069 6411 6103
rect 6561 5117 6595 5151
rect 6377 4981 6411 5015
rect 6193 4777 6227 4811
rect 5273 4709 5307 4743
rect 5489 4709 5523 4743
rect 6469 4709 6503 4743
rect 6009 4641 6043 4675
rect 6285 4641 6319 4675
rect 6377 4641 6411 4675
rect 6561 4641 6595 4675
rect 5641 4505 5675 4539
rect 5457 4437 5491 4471
rect 5825 4437 5859 4471
rect 4997 4165 5031 4199
rect 5917 4029 5951 4063
rect 6193 4029 6227 4063
rect 6561 4029 6595 4063
rect 5457 3961 5491 3995
rect 5825 3961 5859 3995
rect 6377 3893 6411 3927
rect 6101 3689 6135 3723
rect 4905 3621 4939 3655
rect 5273 3621 5307 3655
rect 5917 3621 5951 3655
rect 6285 3621 6319 3655
rect 5089 3553 5123 3587
rect 5365 3553 5399 3587
rect 6193 3553 6227 3587
rect 6469 3485 6503 3519
rect 6377 3145 6411 3179
rect 5917 3009 5951 3043
rect 5365 2941 5399 2975
rect 5457 2941 5491 2975
rect 5641 2941 5675 2975
rect 6193 2941 6227 2975
rect 6561 2941 6595 2975
rect 4813 2873 4847 2907
rect 5273 2601 5307 2635
rect 5441 2601 5475 2635
rect 6193 2601 6227 2635
rect 5641 2533 5675 2567
rect 6009 2465 6043 2499
rect 6285 2465 6319 2499
rect 6561 2465 6595 2499
rect 5917 2397 5951 2431
rect 6101 2397 6135 2431
rect 6377 2329 6411 2363
rect 5457 2261 5491 2295
rect 5273 2057 5307 2091
rect 5365 2057 5399 2091
rect 6377 2057 6411 2091
rect 5089 1853 5123 1887
rect 5273 1853 5307 1887
rect 5549 1853 5583 1887
rect 6009 1853 6043 1887
rect 6193 1853 6227 1887
rect 6561 1853 6595 1887
rect 5733 1785 5767 1819
rect 5825 1785 5859 1819
rect 6377 969 6411 1003
rect 6561 765 6595 799
<< metal1 >>
rect 552 6554 6900 6576
rect 552 6502 3662 6554
rect 3714 6502 3726 6554
rect 3778 6502 3790 6554
rect 3842 6502 3854 6554
rect 3906 6502 3918 6554
rect 3970 6502 6900 6554
rect 552 6480 6900 6502
rect 6270 6196 6276 6248
rect 6328 6196 6334 6248
rect 6546 6196 6552 6248
rect 6604 6196 6610 6248
rect 6086 6060 6092 6112
rect 6144 6060 6150 6112
rect 6365 6103 6423 6109
rect 6365 6069 6377 6103
rect 6411 6100 6423 6103
rect 6638 6100 6644 6112
rect 6411 6072 6644 6100
rect 6411 6069 6423 6072
rect 6365 6063 6423 6069
rect 6638 6060 6644 6072
rect 6696 6060 6702 6112
rect 552 6010 6900 6032
rect 552 5958 4322 6010
rect 4374 5958 4386 6010
rect 4438 5958 4450 6010
rect 4502 5958 4514 6010
rect 4566 5958 4578 6010
rect 4630 5958 6900 6010
rect 552 5936 6900 5958
rect 552 5466 6900 5488
rect 552 5414 3662 5466
rect 3714 5414 3726 5466
rect 3778 5414 3790 5466
rect 3842 5414 3854 5466
rect 3906 5414 3918 5466
rect 3970 5414 6900 5466
rect 552 5392 6900 5414
rect 6546 5108 6552 5160
rect 6604 5108 6610 5160
rect 6362 4972 6368 5024
rect 6420 4972 6426 5024
rect 552 4922 6900 4944
rect 552 4870 4322 4922
rect 4374 4870 4386 4922
rect 4438 4870 4450 4922
rect 4502 4870 4514 4922
rect 4566 4870 4578 4922
rect 4630 4870 6900 4922
rect 552 4848 6900 4870
rect 5902 4808 5908 4820
rect 5276 4780 5908 4808
rect 5276 4749 5304 4780
rect 5902 4768 5908 4780
rect 5960 4808 5966 4820
rect 6086 4808 6092 4820
rect 5960 4780 6092 4808
rect 5960 4768 5966 4780
rect 6086 4768 6092 4780
rect 6144 4808 6150 4820
rect 6181 4811 6239 4817
rect 6181 4808 6193 4811
rect 6144 4780 6193 4808
rect 6144 4768 6150 4780
rect 6181 4777 6193 4780
rect 6227 4777 6239 4811
rect 6181 4771 6239 4777
rect 5261 4743 5319 4749
rect 5261 4709 5273 4743
rect 5307 4709 5319 4743
rect 5261 4703 5319 4709
rect 5477 4743 5535 4749
rect 5477 4709 5489 4743
rect 5523 4740 5535 4743
rect 6457 4743 6515 4749
rect 6457 4740 6469 4743
rect 5523 4712 6132 4740
rect 5523 4709 5535 4712
rect 5477 4703 5535 4709
rect 5997 4675 6055 4681
rect 5997 4641 6009 4675
rect 6043 4641 6055 4675
rect 5997 4635 6055 4641
rect 5629 4539 5687 4545
rect 5629 4505 5641 4539
rect 5675 4536 5687 4539
rect 6012 4536 6040 4635
rect 6104 4616 6132 4712
rect 6288 4712 6469 4740
rect 6288 4681 6316 4712
rect 6457 4709 6469 4712
rect 6503 4709 6515 4743
rect 6457 4703 6515 4709
rect 6273 4675 6331 4681
rect 6273 4641 6285 4675
rect 6319 4641 6331 4675
rect 6273 4635 6331 4641
rect 6362 4632 6368 4684
rect 6420 4632 6426 4684
rect 6549 4675 6607 4681
rect 6549 4641 6561 4675
rect 6595 4672 6607 4675
rect 6638 4672 6644 4684
rect 6595 4644 6644 4672
rect 6595 4641 6607 4644
rect 6549 4635 6607 4641
rect 6638 4632 6644 4644
rect 6696 4632 6702 4684
rect 6086 4564 6092 4616
rect 6144 4604 6150 4616
rect 6380 4604 6408 4632
rect 6144 4576 6408 4604
rect 6144 4564 6150 4576
rect 5675 4508 6040 4536
rect 5675 4505 5687 4508
rect 5629 4499 5687 4505
rect 5445 4471 5503 4477
rect 5445 4437 5457 4471
rect 5491 4468 5503 4471
rect 5534 4468 5540 4480
rect 5491 4440 5540 4468
rect 5491 4437 5503 4440
rect 5445 4431 5503 4437
rect 5534 4428 5540 4440
rect 5592 4428 5598 4480
rect 5810 4428 5816 4480
rect 5868 4428 5874 4480
rect 552 4378 6900 4400
rect 552 4326 3662 4378
rect 3714 4326 3726 4378
rect 3778 4326 3790 4378
rect 3842 4326 3854 4378
rect 3906 4326 3918 4378
rect 3970 4326 6900 4378
rect 552 4304 6900 4326
rect 2774 4156 2780 4208
rect 2832 4196 2838 4208
rect 4985 4199 5043 4205
rect 4985 4196 4997 4199
rect 2832 4168 4997 4196
rect 2832 4156 2838 4168
rect 4985 4165 4997 4168
rect 5031 4165 5043 4199
rect 4985 4159 5043 4165
rect 5902 4020 5908 4072
rect 5960 4020 5966 4072
rect 6178 4020 6184 4072
rect 6236 4020 6242 4072
rect 6546 4020 6552 4072
rect 6604 4020 6610 4072
rect 5074 3952 5080 4004
rect 5132 3992 5138 4004
rect 5445 3995 5503 4001
rect 5445 3992 5457 3995
rect 5132 3964 5457 3992
rect 5132 3952 5138 3964
rect 5445 3961 5457 3964
rect 5491 3961 5503 3995
rect 5445 3955 5503 3961
rect 5534 3952 5540 4004
rect 5592 3992 5598 4004
rect 5813 3995 5871 4001
rect 5813 3992 5825 3995
rect 5592 3964 5825 3992
rect 5592 3952 5598 3964
rect 5813 3961 5825 3964
rect 5859 3992 5871 3995
rect 6270 3992 6276 4004
rect 5859 3964 6276 3992
rect 5859 3961 5871 3964
rect 5813 3955 5871 3961
rect 6270 3952 6276 3964
rect 6328 3992 6334 4004
rect 6638 3992 6644 4004
rect 6328 3964 6644 3992
rect 6328 3952 6334 3964
rect 6638 3952 6644 3964
rect 6696 3952 6702 4004
rect 6362 3884 6368 3936
rect 6420 3884 6426 3936
rect 552 3834 6900 3856
rect 552 3782 4322 3834
rect 4374 3782 4386 3834
rect 4438 3782 4450 3834
rect 4502 3782 4514 3834
rect 4566 3782 4578 3834
rect 4630 3782 6900 3834
rect 552 3760 6900 3782
rect 5994 3680 6000 3732
rect 6052 3720 6058 3732
rect 6089 3723 6147 3729
rect 6089 3720 6101 3723
rect 6052 3692 6101 3720
rect 6052 3680 6058 3692
rect 6089 3689 6101 3692
rect 6135 3720 6147 3723
rect 6362 3720 6368 3732
rect 6135 3692 6368 3720
rect 6135 3689 6147 3692
rect 6089 3683 6147 3689
rect 6362 3680 6368 3692
rect 6420 3680 6426 3732
rect 4154 3612 4160 3664
rect 4212 3652 4218 3664
rect 4893 3655 4951 3661
rect 4893 3652 4905 3655
rect 4212 3624 4905 3652
rect 4212 3612 4218 3624
rect 4893 3621 4905 3624
rect 4939 3621 4951 3655
rect 4893 3615 4951 3621
rect 5261 3655 5319 3661
rect 5261 3621 5273 3655
rect 5307 3652 5319 3655
rect 5442 3652 5448 3664
rect 5307 3624 5448 3652
rect 5307 3621 5319 3624
rect 5261 3615 5319 3621
rect 5442 3612 5448 3624
rect 5500 3652 5506 3664
rect 5905 3655 5963 3661
rect 5905 3652 5917 3655
rect 5500 3624 5917 3652
rect 5500 3612 5506 3624
rect 5905 3621 5917 3624
rect 5951 3621 5963 3655
rect 5905 3615 5963 3621
rect 6270 3612 6276 3664
rect 6328 3612 6334 3664
rect 5074 3544 5080 3596
rect 5132 3544 5138 3596
rect 5353 3587 5411 3593
rect 5353 3553 5365 3587
rect 5399 3553 5411 3587
rect 5353 3547 5411 3553
rect 5258 3476 5264 3528
rect 5316 3516 5322 3528
rect 5368 3516 5396 3547
rect 6086 3544 6092 3596
rect 6144 3584 6150 3596
rect 6181 3587 6239 3593
rect 6181 3584 6193 3587
rect 6144 3556 6193 3584
rect 6144 3544 6150 3556
rect 6181 3553 6193 3556
rect 6227 3553 6239 3587
rect 6181 3547 6239 3553
rect 5316 3488 5396 3516
rect 5316 3476 5322 3488
rect 5902 3476 5908 3528
rect 5960 3516 5966 3528
rect 6457 3519 6515 3525
rect 6457 3516 6469 3519
rect 5960 3488 6469 3516
rect 5960 3476 5966 3488
rect 6457 3485 6469 3488
rect 6503 3485 6515 3519
rect 6457 3479 6515 3485
rect 552 3290 6900 3312
rect 552 3238 3662 3290
rect 3714 3238 3726 3290
rect 3778 3238 3790 3290
rect 3842 3238 3854 3290
rect 3906 3238 3918 3290
rect 3970 3238 6900 3290
rect 552 3216 6900 3238
rect 6178 3136 6184 3188
rect 6236 3176 6242 3188
rect 6365 3179 6423 3185
rect 6365 3176 6377 3179
rect 6236 3148 6377 3176
rect 6236 3136 6242 3148
rect 6365 3145 6377 3148
rect 6411 3145 6423 3179
rect 6365 3139 6423 3145
rect 5810 3000 5816 3052
rect 5868 3040 5874 3052
rect 5905 3043 5963 3049
rect 5905 3040 5917 3043
rect 5868 3012 5917 3040
rect 5868 3000 5874 3012
rect 5905 3009 5917 3012
rect 5951 3009 5963 3043
rect 5905 3003 5963 3009
rect 5350 2932 5356 2984
rect 5408 2932 5414 2984
rect 5442 2932 5448 2984
rect 5500 2932 5506 2984
rect 5626 2932 5632 2984
rect 5684 2932 5690 2984
rect 6178 2932 6184 2984
rect 6236 2972 6242 2984
rect 6549 2975 6607 2981
rect 6549 2972 6561 2975
rect 6236 2944 6561 2972
rect 6236 2932 6242 2944
rect 6549 2941 6561 2944
rect 6595 2941 6607 2975
rect 6549 2935 6607 2941
rect 4798 2864 4804 2916
rect 4856 2864 4862 2916
rect 552 2746 6900 2768
rect 552 2694 4322 2746
rect 4374 2694 4386 2746
rect 4438 2694 4450 2746
rect 4502 2694 4514 2746
rect 4566 2694 4578 2746
rect 4630 2694 6900 2746
rect 552 2672 6900 2694
rect 5074 2592 5080 2644
rect 5132 2632 5138 2644
rect 5442 2641 5448 2644
rect 5261 2635 5319 2641
rect 5261 2632 5273 2635
rect 5132 2604 5273 2632
rect 5132 2592 5138 2604
rect 5261 2601 5273 2604
rect 5307 2601 5319 2635
rect 5261 2595 5319 2601
rect 5429 2635 5448 2641
rect 5429 2601 5441 2635
rect 5429 2595 5448 2601
rect 5442 2592 5448 2595
rect 5500 2592 5506 2644
rect 6178 2592 6184 2644
rect 6236 2592 6242 2644
rect 5626 2524 5632 2576
rect 5684 2564 5690 2576
rect 5684 2536 6132 2564
rect 5684 2524 5690 2536
rect 5994 2456 6000 2508
rect 6052 2456 6058 2508
rect 6104 2437 6132 2536
rect 6273 2499 6331 2505
rect 6273 2465 6285 2499
rect 6319 2496 6331 2499
rect 6362 2496 6368 2508
rect 6319 2468 6368 2496
rect 6319 2465 6331 2468
rect 6273 2459 6331 2465
rect 6362 2456 6368 2468
rect 6420 2456 6426 2508
rect 6546 2456 6552 2508
rect 6604 2456 6610 2508
rect 5905 2431 5963 2437
rect 5905 2397 5917 2431
rect 5951 2397 5963 2431
rect 5905 2391 5963 2397
rect 6089 2431 6147 2437
rect 6089 2397 6101 2431
rect 6135 2428 6147 2431
rect 6135 2400 6408 2428
rect 6135 2397 6147 2400
rect 6089 2391 6147 2397
rect 5920 2360 5948 2391
rect 6178 2360 6184 2372
rect 5920 2332 6184 2360
rect 6178 2320 6184 2332
rect 6236 2320 6242 2372
rect 6380 2369 6408 2400
rect 6365 2363 6423 2369
rect 6365 2329 6377 2363
rect 6411 2329 6423 2363
rect 6365 2323 6423 2329
rect 5445 2295 5503 2301
rect 5445 2261 5457 2295
rect 5491 2292 5503 2295
rect 6270 2292 6276 2304
rect 5491 2264 6276 2292
rect 5491 2261 5503 2264
rect 5445 2255 5503 2261
rect 6270 2252 6276 2264
rect 6328 2252 6334 2304
rect 552 2202 6900 2224
rect 552 2150 3662 2202
rect 3714 2150 3726 2202
rect 3778 2150 3790 2202
rect 3842 2150 3854 2202
rect 3906 2150 3918 2202
rect 3970 2150 6900 2202
rect 552 2128 6900 2150
rect 5258 2048 5264 2100
rect 5316 2048 5322 2100
rect 5350 2048 5356 2100
rect 5408 2048 5414 2100
rect 6362 2048 6368 2100
rect 6420 2048 6426 2100
rect 5276 1952 5304 2048
rect 6380 1952 6408 2048
rect 5276 1924 5580 1952
rect 5552 1893 5580 1924
rect 6012 1924 6408 1952
rect 6012 1893 6040 1924
rect 5077 1887 5135 1893
rect 5077 1853 5089 1887
rect 5123 1853 5135 1887
rect 5077 1847 5135 1853
rect 5261 1887 5319 1893
rect 5261 1853 5273 1887
rect 5307 1853 5319 1887
rect 5261 1847 5319 1853
rect 5537 1887 5595 1893
rect 5537 1853 5549 1887
rect 5583 1853 5595 1887
rect 5997 1887 6055 1893
rect 5997 1884 6009 1887
rect 5537 1847 5595 1853
rect 5644 1856 6009 1884
rect 5092 1748 5120 1847
rect 5276 1816 5304 1847
rect 5644 1816 5672 1856
rect 5997 1853 6009 1856
rect 6043 1853 6055 1887
rect 5997 1847 6055 1853
rect 6178 1844 6184 1896
rect 6236 1884 6242 1896
rect 6362 1884 6368 1896
rect 6236 1856 6368 1884
rect 6236 1844 6242 1856
rect 6362 1844 6368 1856
rect 6420 1844 6426 1896
rect 6546 1844 6552 1896
rect 6604 1844 6610 1896
rect 5276 1788 5672 1816
rect 5721 1819 5779 1825
rect 5721 1785 5733 1819
rect 5767 1816 5779 1819
rect 5813 1819 5871 1825
rect 5813 1816 5825 1819
rect 5767 1788 5825 1816
rect 5767 1785 5779 1788
rect 5721 1779 5779 1785
rect 5813 1785 5825 1788
rect 5859 1785 5871 1819
rect 5813 1779 5871 1785
rect 6196 1748 6224 1844
rect 5092 1720 6224 1748
rect 552 1658 6900 1680
rect 552 1606 4322 1658
rect 4374 1606 4386 1658
rect 4438 1606 4450 1658
rect 4502 1606 4514 1658
rect 4566 1606 4578 1658
rect 4630 1606 6900 1658
rect 552 1584 6900 1606
rect 552 1114 6900 1136
rect 552 1062 3662 1114
rect 3714 1062 3726 1114
rect 3778 1062 3790 1114
rect 3842 1062 3854 1114
rect 3906 1062 3918 1114
rect 3970 1062 6900 1114
rect 552 1040 6900 1062
rect 6362 960 6368 1012
rect 6420 960 6426 1012
rect 6546 756 6552 808
rect 6604 756 6610 808
rect 552 570 6900 592
rect 552 518 4322 570
rect 4374 518 4386 570
rect 4438 518 4450 570
rect 4502 518 4514 570
rect 4566 518 4578 570
rect 4630 518 6900 570
rect 552 496 6900 518
<< via1 >>
rect 3662 6502 3714 6554
rect 3726 6502 3778 6554
rect 3790 6502 3842 6554
rect 3854 6502 3906 6554
rect 3918 6502 3970 6554
rect 6276 6239 6328 6248
rect 6276 6205 6285 6239
rect 6285 6205 6319 6239
rect 6319 6205 6328 6239
rect 6276 6196 6328 6205
rect 6552 6239 6604 6248
rect 6552 6205 6561 6239
rect 6561 6205 6595 6239
rect 6595 6205 6604 6239
rect 6552 6196 6604 6205
rect 6092 6103 6144 6112
rect 6092 6069 6101 6103
rect 6101 6069 6135 6103
rect 6135 6069 6144 6103
rect 6092 6060 6144 6069
rect 6644 6060 6696 6112
rect 4322 5958 4374 6010
rect 4386 5958 4438 6010
rect 4450 5958 4502 6010
rect 4514 5958 4566 6010
rect 4578 5958 4630 6010
rect 3662 5414 3714 5466
rect 3726 5414 3778 5466
rect 3790 5414 3842 5466
rect 3854 5414 3906 5466
rect 3918 5414 3970 5466
rect 6552 5151 6604 5160
rect 6552 5117 6561 5151
rect 6561 5117 6595 5151
rect 6595 5117 6604 5151
rect 6552 5108 6604 5117
rect 6368 5015 6420 5024
rect 6368 4981 6377 5015
rect 6377 4981 6411 5015
rect 6411 4981 6420 5015
rect 6368 4972 6420 4981
rect 4322 4870 4374 4922
rect 4386 4870 4438 4922
rect 4450 4870 4502 4922
rect 4514 4870 4566 4922
rect 4578 4870 4630 4922
rect 5908 4768 5960 4820
rect 6092 4768 6144 4820
rect 6368 4675 6420 4684
rect 6368 4641 6377 4675
rect 6377 4641 6411 4675
rect 6411 4641 6420 4675
rect 6368 4632 6420 4641
rect 6644 4632 6696 4684
rect 6092 4564 6144 4616
rect 5540 4428 5592 4480
rect 5816 4471 5868 4480
rect 5816 4437 5825 4471
rect 5825 4437 5859 4471
rect 5859 4437 5868 4471
rect 5816 4428 5868 4437
rect 3662 4326 3714 4378
rect 3726 4326 3778 4378
rect 3790 4326 3842 4378
rect 3854 4326 3906 4378
rect 3918 4326 3970 4378
rect 2780 4156 2832 4208
rect 5908 4063 5960 4072
rect 5908 4029 5917 4063
rect 5917 4029 5951 4063
rect 5951 4029 5960 4063
rect 5908 4020 5960 4029
rect 6184 4063 6236 4072
rect 6184 4029 6193 4063
rect 6193 4029 6227 4063
rect 6227 4029 6236 4063
rect 6184 4020 6236 4029
rect 6552 4063 6604 4072
rect 6552 4029 6561 4063
rect 6561 4029 6595 4063
rect 6595 4029 6604 4063
rect 6552 4020 6604 4029
rect 5080 3952 5132 4004
rect 5540 3952 5592 4004
rect 6276 3952 6328 4004
rect 6644 3952 6696 4004
rect 6368 3927 6420 3936
rect 6368 3893 6377 3927
rect 6377 3893 6411 3927
rect 6411 3893 6420 3927
rect 6368 3884 6420 3893
rect 4322 3782 4374 3834
rect 4386 3782 4438 3834
rect 4450 3782 4502 3834
rect 4514 3782 4566 3834
rect 4578 3782 4630 3834
rect 6000 3680 6052 3732
rect 6368 3680 6420 3732
rect 4160 3612 4212 3664
rect 5448 3612 5500 3664
rect 6276 3655 6328 3664
rect 6276 3621 6285 3655
rect 6285 3621 6319 3655
rect 6319 3621 6328 3655
rect 6276 3612 6328 3621
rect 5080 3587 5132 3596
rect 5080 3553 5089 3587
rect 5089 3553 5123 3587
rect 5123 3553 5132 3587
rect 5080 3544 5132 3553
rect 5264 3476 5316 3528
rect 6092 3544 6144 3596
rect 5908 3476 5960 3528
rect 3662 3238 3714 3290
rect 3726 3238 3778 3290
rect 3790 3238 3842 3290
rect 3854 3238 3906 3290
rect 3918 3238 3970 3290
rect 6184 3136 6236 3188
rect 5816 3000 5868 3052
rect 5356 2975 5408 2984
rect 5356 2941 5365 2975
rect 5365 2941 5399 2975
rect 5399 2941 5408 2975
rect 5356 2932 5408 2941
rect 5448 2975 5500 2984
rect 5448 2941 5457 2975
rect 5457 2941 5491 2975
rect 5491 2941 5500 2975
rect 5448 2932 5500 2941
rect 5632 2975 5684 2984
rect 5632 2941 5641 2975
rect 5641 2941 5675 2975
rect 5675 2941 5684 2975
rect 5632 2932 5684 2941
rect 6184 2975 6236 2984
rect 6184 2941 6193 2975
rect 6193 2941 6227 2975
rect 6227 2941 6236 2975
rect 6184 2932 6236 2941
rect 4804 2907 4856 2916
rect 4804 2873 4813 2907
rect 4813 2873 4847 2907
rect 4847 2873 4856 2907
rect 4804 2864 4856 2873
rect 4322 2694 4374 2746
rect 4386 2694 4438 2746
rect 4450 2694 4502 2746
rect 4514 2694 4566 2746
rect 4578 2694 4630 2746
rect 5080 2592 5132 2644
rect 5448 2635 5500 2644
rect 5448 2601 5475 2635
rect 5475 2601 5500 2635
rect 5448 2592 5500 2601
rect 6184 2635 6236 2644
rect 6184 2601 6193 2635
rect 6193 2601 6227 2635
rect 6227 2601 6236 2635
rect 6184 2592 6236 2601
rect 5632 2567 5684 2576
rect 5632 2533 5641 2567
rect 5641 2533 5675 2567
rect 5675 2533 5684 2567
rect 5632 2524 5684 2533
rect 6000 2499 6052 2508
rect 6000 2465 6009 2499
rect 6009 2465 6043 2499
rect 6043 2465 6052 2499
rect 6000 2456 6052 2465
rect 6368 2456 6420 2508
rect 6552 2499 6604 2508
rect 6552 2465 6561 2499
rect 6561 2465 6595 2499
rect 6595 2465 6604 2499
rect 6552 2456 6604 2465
rect 6184 2320 6236 2372
rect 6276 2252 6328 2304
rect 3662 2150 3714 2202
rect 3726 2150 3778 2202
rect 3790 2150 3842 2202
rect 3854 2150 3906 2202
rect 3918 2150 3970 2202
rect 5264 2091 5316 2100
rect 5264 2057 5273 2091
rect 5273 2057 5307 2091
rect 5307 2057 5316 2091
rect 5264 2048 5316 2057
rect 5356 2091 5408 2100
rect 5356 2057 5365 2091
rect 5365 2057 5399 2091
rect 5399 2057 5408 2091
rect 5356 2048 5408 2057
rect 6368 2091 6420 2100
rect 6368 2057 6377 2091
rect 6377 2057 6411 2091
rect 6411 2057 6420 2091
rect 6368 2048 6420 2057
rect 6184 1887 6236 1896
rect 6184 1853 6193 1887
rect 6193 1853 6227 1887
rect 6227 1853 6236 1887
rect 6184 1844 6236 1853
rect 6368 1844 6420 1896
rect 6552 1887 6604 1896
rect 6552 1853 6561 1887
rect 6561 1853 6595 1887
rect 6595 1853 6604 1887
rect 6552 1844 6604 1853
rect 4322 1606 4374 1658
rect 4386 1606 4438 1658
rect 4450 1606 4502 1658
rect 4514 1606 4566 1658
rect 4578 1606 4630 1658
rect 3662 1062 3714 1114
rect 3726 1062 3778 1114
rect 3790 1062 3842 1114
rect 3854 1062 3906 1114
rect 3918 1062 3970 1114
rect 6368 1003 6420 1012
rect 6368 969 6377 1003
rect 6377 969 6411 1003
rect 6411 969 6420 1003
rect 6368 960 6420 969
rect 6552 799 6604 808
rect 6552 765 6561 799
rect 6561 765 6595 799
rect 6595 765 6604 799
rect 6552 756 6604 765
rect 4322 518 4374 570
rect 4386 518 4438 570
rect 4450 518 4502 570
rect 4514 518 4566 570
rect 4578 518 4630 570
<< metal2 >>
rect 6274 6624 6330 6633
rect 3662 6556 3970 6565
rect 6274 6559 6330 6568
rect 3662 6554 3668 6556
rect 3724 6554 3748 6556
rect 3804 6554 3828 6556
rect 3884 6554 3908 6556
rect 3964 6554 3970 6556
rect 3724 6502 3726 6554
rect 3906 6502 3908 6554
rect 3662 6500 3668 6502
rect 3724 6500 3748 6502
rect 3804 6500 3828 6502
rect 3884 6500 3908 6502
rect 3964 6500 3970 6502
rect 3662 6491 3970 6500
rect 6288 6254 6316 6559
rect 6276 6248 6328 6254
rect 6276 6190 6328 6196
rect 6552 6248 6604 6254
rect 6552 6190 6604 6196
rect 6092 6112 6144 6118
rect 4158 6080 4214 6089
rect 6564 6089 6592 6190
rect 6644 6112 6696 6118
rect 6092 6054 6144 6060
rect 6550 6080 6606 6089
rect 4158 6015 4214 6024
rect 3662 5468 3970 5477
rect 3662 5466 3668 5468
rect 3724 5466 3748 5468
rect 3804 5466 3828 5468
rect 3884 5466 3908 5468
rect 3964 5466 3970 5468
rect 3724 5414 3726 5466
rect 3906 5414 3908 5466
rect 3662 5412 3668 5414
rect 3724 5412 3748 5414
rect 3804 5412 3828 5414
rect 3884 5412 3908 5414
rect 3964 5412 3970 5414
rect 3662 5403 3970 5412
rect 3662 4380 3970 4389
rect 3662 4378 3668 4380
rect 3724 4378 3748 4380
rect 3804 4378 3828 4380
rect 3884 4378 3908 4380
rect 3964 4378 3970 4380
rect 3724 4326 3726 4378
rect 3906 4326 3908 4378
rect 3662 4324 3668 4326
rect 3724 4324 3748 4326
rect 3804 4324 3828 4326
rect 3884 4324 3908 4326
rect 3964 4324 3970 4326
rect 3662 4315 3970 4324
rect 2780 4208 2832 4214
rect 2780 4150 2832 4156
rect 2792 3641 2820 4150
rect 4172 3670 4200 6015
rect 4322 6012 4630 6021
rect 4322 6010 4328 6012
rect 4384 6010 4408 6012
rect 4464 6010 4488 6012
rect 4544 6010 4568 6012
rect 4624 6010 4630 6012
rect 4384 5958 4386 6010
rect 4566 5958 4568 6010
rect 4322 5956 4328 5958
rect 4384 5956 4408 5958
rect 4464 5956 4488 5958
rect 4544 5956 4568 5958
rect 4624 5956 4630 5958
rect 4322 5947 4630 5956
rect 4322 4924 4630 4933
rect 4322 4922 4328 4924
rect 4384 4922 4408 4924
rect 4464 4922 4488 4924
rect 4544 4922 4568 4924
rect 4624 4922 4630 4924
rect 4384 4870 4386 4922
rect 4566 4870 4568 4922
rect 4322 4868 4328 4870
rect 4384 4868 4408 4870
rect 4464 4868 4488 4870
rect 4544 4868 4568 4870
rect 4624 4868 4630 4870
rect 4322 4859 4630 4868
rect 6104 4826 6132 6054
rect 6644 6054 6696 6060
rect 6550 6015 6606 6024
rect 6552 5160 6604 5166
rect 6552 5102 6604 5108
rect 6368 5024 6420 5030
rect 6564 5001 6592 5102
rect 6368 4966 6420 4972
rect 6550 4992 6606 5001
rect 5908 4820 5960 4826
rect 5908 4762 5960 4768
rect 6092 4820 6144 4826
rect 6092 4762 6144 4768
rect 5540 4480 5592 4486
rect 5540 4422 5592 4428
rect 5816 4480 5868 4486
rect 5816 4422 5868 4428
rect 5552 4010 5580 4422
rect 5080 4004 5132 4010
rect 5080 3946 5132 3952
rect 5540 4004 5592 4010
rect 5540 3946 5592 3952
rect 4322 3836 4630 3845
rect 4322 3834 4328 3836
rect 4384 3834 4408 3836
rect 4464 3834 4488 3836
rect 4544 3834 4568 3836
rect 4624 3834 4630 3836
rect 4384 3782 4386 3834
rect 4566 3782 4568 3834
rect 4322 3780 4328 3782
rect 4384 3780 4408 3782
rect 4464 3780 4488 3782
rect 4544 3780 4568 3782
rect 4624 3780 4630 3782
rect 4322 3771 4630 3780
rect 4160 3664 4212 3670
rect 2778 3632 2834 3641
rect 4160 3606 4212 3612
rect 5092 3602 5120 3946
rect 5448 3664 5500 3670
rect 5448 3606 5500 3612
rect 2778 3567 2834 3576
rect 5080 3596 5132 3602
rect 5080 3538 5132 3544
rect 3662 3292 3970 3301
rect 3662 3290 3668 3292
rect 3724 3290 3748 3292
rect 3804 3290 3828 3292
rect 3884 3290 3908 3292
rect 3964 3290 3970 3292
rect 3724 3238 3726 3290
rect 3906 3238 3908 3290
rect 3662 3236 3668 3238
rect 3724 3236 3748 3238
rect 3804 3236 3828 3238
rect 3884 3236 3908 3238
rect 3964 3236 3970 3238
rect 3662 3227 3970 3236
rect 4804 2916 4856 2922
rect 4804 2858 4856 2864
rect 4322 2748 4630 2757
rect 4322 2746 4328 2748
rect 4384 2746 4408 2748
rect 4464 2746 4488 2748
rect 4544 2746 4568 2748
rect 4624 2746 4630 2748
rect 4384 2694 4386 2746
rect 4566 2694 4568 2746
rect 4322 2692 4328 2694
rect 4384 2692 4408 2694
rect 4464 2692 4488 2694
rect 4544 2692 4568 2694
rect 4624 2692 4630 2694
rect 4322 2683 4630 2692
rect 3662 2204 3970 2213
rect 3662 2202 3668 2204
rect 3724 2202 3748 2204
rect 3804 2202 3828 2204
rect 3884 2202 3908 2204
rect 3964 2202 3970 2204
rect 3724 2150 3726 2202
rect 3906 2150 3908 2202
rect 3662 2148 3668 2150
rect 3724 2148 3748 2150
rect 3804 2148 3828 2150
rect 3884 2148 3908 2150
rect 3964 2148 3970 2150
rect 3662 2139 3970 2148
rect 4322 1660 4630 1669
rect 4322 1658 4328 1660
rect 4384 1658 4408 1660
rect 4464 1658 4488 1660
rect 4544 1658 4568 1660
rect 4624 1658 4630 1660
rect 4384 1606 4386 1658
rect 4566 1606 4568 1658
rect 4322 1604 4328 1606
rect 4384 1604 4408 1606
rect 4464 1604 4488 1606
rect 4544 1604 4568 1606
rect 4624 1604 4630 1606
rect 4322 1595 4630 1604
rect 4816 1329 4844 2858
rect 5092 2650 5120 3538
rect 5264 3528 5316 3534
rect 5264 3470 5316 3476
rect 5080 2644 5132 2650
rect 5080 2586 5132 2592
rect 5276 2106 5304 3470
rect 5460 2990 5488 3606
rect 5828 3058 5856 4422
rect 5920 4078 5948 4762
rect 6380 4690 6408 4966
rect 6550 4927 6606 4936
rect 6656 4690 6684 6054
rect 6368 4684 6420 4690
rect 6368 4626 6420 4632
rect 6644 4684 6696 4690
rect 6644 4626 6696 4632
rect 6092 4616 6144 4622
rect 6092 4558 6144 4564
rect 5908 4072 5960 4078
rect 5908 4014 5960 4020
rect 5920 3534 5948 4014
rect 6000 3732 6052 3738
rect 6000 3674 6052 3680
rect 5908 3528 5960 3534
rect 5908 3470 5960 3476
rect 5816 3052 5868 3058
rect 5816 2994 5868 3000
rect 5356 2984 5408 2990
rect 5356 2926 5408 2932
rect 5448 2984 5500 2990
rect 5448 2926 5500 2932
rect 5632 2984 5684 2990
rect 5632 2926 5684 2932
rect 5368 2106 5396 2926
rect 5460 2650 5488 2926
rect 5448 2644 5500 2650
rect 5448 2586 5500 2592
rect 5644 2582 5672 2926
rect 5632 2576 5684 2582
rect 5632 2518 5684 2524
rect 6012 2514 6040 3674
rect 6104 3602 6132 4558
rect 6184 4072 6236 4078
rect 6184 4014 6236 4020
rect 6552 4072 6604 4078
rect 6552 4014 6604 4020
rect 6092 3596 6144 3602
rect 6092 3538 6144 3544
rect 6196 3194 6224 4014
rect 6276 4004 6328 4010
rect 6276 3946 6328 3952
rect 6288 3670 6316 3946
rect 6368 3936 6420 3942
rect 6564 3913 6592 4014
rect 6656 4010 6684 4626
rect 6644 4004 6696 4010
rect 6644 3946 6696 3952
rect 6368 3878 6420 3884
rect 6550 3904 6606 3913
rect 6380 3738 6408 3878
rect 6550 3839 6606 3848
rect 6368 3732 6420 3738
rect 6368 3674 6420 3680
rect 6276 3664 6328 3670
rect 6276 3606 6328 3612
rect 6184 3188 6236 3194
rect 6184 3130 6236 3136
rect 6184 2984 6236 2990
rect 6184 2926 6236 2932
rect 6196 2650 6224 2926
rect 6184 2644 6236 2650
rect 6184 2586 6236 2592
rect 6550 2544 6606 2553
rect 6000 2508 6052 2514
rect 6000 2450 6052 2456
rect 6368 2508 6420 2514
rect 6550 2479 6552 2488
rect 6368 2450 6420 2456
rect 6604 2479 6606 2488
rect 6552 2450 6604 2456
rect 6184 2372 6236 2378
rect 6184 2314 6236 2320
rect 5264 2100 5316 2106
rect 5264 2042 5316 2048
rect 5356 2100 5408 2106
rect 5356 2042 5408 2048
rect 6196 1902 6224 2314
rect 6276 2304 6328 2310
rect 6380 2258 6408 2450
rect 6328 2252 6408 2258
rect 6276 2246 6408 2252
rect 6288 2230 6408 2246
rect 6380 2106 6408 2230
rect 6368 2100 6420 2106
rect 6368 2042 6420 2048
rect 6184 1896 6236 1902
rect 6184 1838 6236 1844
rect 6368 1896 6420 1902
rect 6368 1838 6420 1844
rect 6552 1896 6604 1902
rect 6552 1838 6604 1844
rect 4802 1320 4858 1329
rect 4802 1255 4858 1264
rect 3662 1116 3970 1125
rect 3662 1114 3668 1116
rect 3724 1114 3748 1116
rect 3804 1114 3828 1116
rect 3884 1114 3908 1116
rect 3964 1114 3970 1116
rect 3724 1062 3726 1114
rect 3906 1062 3908 1114
rect 3662 1060 3668 1062
rect 3724 1060 3748 1062
rect 3804 1060 3828 1062
rect 3884 1060 3908 1062
rect 3964 1060 3970 1062
rect 3662 1051 3970 1060
rect 6380 1018 6408 1838
rect 6564 1737 6592 1838
rect 6550 1728 6606 1737
rect 6550 1663 6606 1672
rect 6368 1012 6420 1018
rect 6368 954 6420 960
rect 6552 808 6604 814
rect 6552 750 6604 756
rect 6564 649 6592 750
rect 6550 640 6606 649
rect 4322 572 4630 581
rect 6550 575 6606 584
rect 4322 570 4328 572
rect 4384 570 4408 572
rect 4464 570 4488 572
rect 4544 570 4568 572
rect 4624 570 4630 572
rect 4384 518 4386 570
rect 4566 518 4568 570
rect 4322 516 4328 518
rect 4384 516 4408 518
rect 4464 516 4488 518
rect 4544 516 4568 518
rect 4624 516 4630 518
rect 4322 507 4630 516
rect 3698 0 3754 400
<< via2 >>
rect 6274 6568 6330 6624
rect 3668 6554 3724 6556
rect 3748 6554 3804 6556
rect 3828 6554 3884 6556
rect 3908 6554 3964 6556
rect 3668 6502 3714 6554
rect 3714 6502 3724 6554
rect 3748 6502 3778 6554
rect 3778 6502 3790 6554
rect 3790 6502 3804 6554
rect 3828 6502 3842 6554
rect 3842 6502 3854 6554
rect 3854 6502 3884 6554
rect 3908 6502 3918 6554
rect 3918 6502 3964 6554
rect 3668 6500 3724 6502
rect 3748 6500 3804 6502
rect 3828 6500 3884 6502
rect 3908 6500 3964 6502
rect 4158 6024 4214 6080
rect 3668 5466 3724 5468
rect 3748 5466 3804 5468
rect 3828 5466 3884 5468
rect 3908 5466 3964 5468
rect 3668 5414 3714 5466
rect 3714 5414 3724 5466
rect 3748 5414 3778 5466
rect 3778 5414 3790 5466
rect 3790 5414 3804 5466
rect 3828 5414 3842 5466
rect 3842 5414 3854 5466
rect 3854 5414 3884 5466
rect 3908 5414 3918 5466
rect 3918 5414 3964 5466
rect 3668 5412 3724 5414
rect 3748 5412 3804 5414
rect 3828 5412 3884 5414
rect 3908 5412 3964 5414
rect 3668 4378 3724 4380
rect 3748 4378 3804 4380
rect 3828 4378 3884 4380
rect 3908 4378 3964 4380
rect 3668 4326 3714 4378
rect 3714 4326 3724 4378
rect 3748 4326 3778 4378
rect 3778 4326 3790 4378
rect 3790 4326 3804 4378
rect 3828 4326 3842 4378
rect 3842 4326 3854 4378
rect 3854 4326 3884 4378
rect 3908 4326 3918 4378
rect 3918 4326 3964 4378
rect 3668 4324 3724 4326
rect 3748 4324 3804 4326
rect 3828 4324 3884 4326
rect 3908 4324 3964 4326
rect 4328 6010 4384 6012
rect 4408 6010 4464 6012
rect 4488 6010 4544 6012
rect 4568 6010 4624 6012
rect 4328 5958 4374 6010
rect 4374 5958 4384 6010
rect 4408 5958 4438 6010
rect 4438 5958 4450 6010
rect 4450 5958 4464 6010
rect 4488 5958 4502 6010
rect 4502 5958 4514 6010
rect 4514 5958 4544 6010
rect 4568 5958 4578 6010
rect 4578 5958 4624 6010
rect 4328 5956 4384 5958
rect 4408 5956 4464 5958
rect 4488 5956 4544 5958
rect 4568 5956 4624 5958
rect 4328 4922 4384 4924
rect 4408 4922 4464 4924
rect 4488 4922 4544 4924
rect 4568 4922 4624 4924
rect 4328 4870 4374 4922
rect 4374 4870 4384 4922
rect 4408 4870 4438 4922
rect 4438 4870 4450 4922
rect 4450 4870 4464 4922
rect 4488 4870 4502 4922
rect 4502 4870 4514 4922
rect 4514 4870 4544 4922
rect 4568 4870 4578 4922
rect 4578 4870 4624 4922
rect 4328 4868 4384 4870
rect 4408 4868 4464 4870
rect 4488 4868 4544 4870
rect 4568 4868 4624 4870
rect 6550 6024 6606 6080
rect 4328 3834 4384 3836
rect 4408 3834 4464 3836
rect 4488 3834 4544 3836
rect 4568 3834 4624 3836
rect 4328 3782 4374 3834
rect 4374 3782 4384 3834
rect 4408 3782 4438 3834
rect 4438 3782 4450 3834
rect 4450 3782 4464 3834
rect 4488 3782 4502 3834
rect 4502 3782 4514 3834
rect 4514 3782 4544 3834
rect 4568 3782 4578 3834
rect 4578 3782 4624 3834
rect 4328 3780 4384 3782
rect 4408 3780 4464 3782
rect 4488 3780 4544 3782
rect 4568 3780 4624 3782
rect 2778 3576 2834 3632
rect 3668 3290 3724 3292
rect 3748 3290 3804 3292
rect 3828 3290 3884 3292
rect 3908 3290 3964 3292
rect 3668 3238 3714 3290
rect 3714 3238 3724 3290
rect 3748 3238 3778 3290
rect 3778 3238 3790 3290
rect 3790 3238 3804 3290
rect 3828 3238 3842 3290
rect 3842 3238 3854 3290
rect 3854 3238 3884 3290
rect 3908 3238 3918 3290
rect 3918 3238 3964 3290
rect 3668 3236 3724 3238
rect 3748 3236 3804 3238
rect 3828 3236 3884 3238
rect 3908 3236 3964 3238
rect 4328 2746 4384 2748
rect 4408 2746 4464 2748
rect 4488 2746 4544 2748
rect 4568 2746 4624 2748
rect 4328 2694 4374 2746
rect 4374 2694 4384 2746
rect 4408 2694 4438 2746
rect 4438 2694 4450 2746
rect 4450 2694 4464 2746
rect 4488 2694 4502 2746
rect 4502 2694 4514 2746
rect 4514 2694 4544 2746
rect 4568 2694 4578 2746
rect 4578 2694 4624 2746
rect 4328 2692 4384 2694
rect 4408 2692 4464 2694
rect 4488 2692 4544 2694
rect 4568 2692 4624 2694
rect 3668 2202 3724 2204
rect 3748 2202 3804 2204
rect 3828 2202 3884 2204
rect 3908 2202 3964 2204
rect 3668 2150 3714 2202
rect 3714 2150 3724 2202
rect 3748 2150 3778 2202
rect 3778 2150 3790 2202
rect 3790 2150 3804 2202
rect 3828 2150 3842 2202
rect 3842 2150 3854 2202
rect 3854 2150 3884 2202
rect 3908 2150 3918 2202
rect 3918 2150 3964 2202
rect 3668 2148 3724 2150
rect 3748 2148 3804 2150
rect 3828 2148 3884 2150
rect 3908 2148 3964 2150
rect 4328 1658 4384 1660
rect 4408 1658 4464 1660
rect 4488 1658 4544 1660
rect 4568 1658 4624 1660
rect 4328 1606 4374 1658
rect 4374 1606 4384 1658
rect 4408 1606 4438 1658
rect 4438 1606 4450 1658
rect 4450 1606 4464 1658
rect 4488 1606 4502 1658
rect 4502 1606 4514 1658
rect 4514 1606 4544 1658
rect 4568 1606 4578 1658
rect 4578 1606 4624 1658
rect 4328 1604 4384 1606
rect 4408 1604 4464 1606
rect 4488 1604 4544 1606
rect 4568 1604 4624 1606
rect 6550 4936 6606 4992
rect 6550 3848 6606 3904
rect 6550 2508 6606 2544
rect 6550 2488 6552 2508
rect 6552 2488 6604 2508
rect 6604 2488 6606 2508
rect 4802 1264 4858 1320
rect 3668 1114 3724 1116
rect 3748 1114 3804 1116
rect 3828 1114 3884 1116
rect 3908 1114 3964 1116
rect 3668 1062 3714 1114
rect 3714 1062 3724 1114
rect 3748 1062 3778 1114
rect 3778 1062 3790 1114
rect 3790 1062 3804 1114
rect 3828 1062 3842 1114
rect 3842 1062 3854 1114
rect 3854 1062 3884 1114
rect 3908 1062 3918 1114
rect 3918 1062 3964 1114
rect 3668 1060 3724 1062
rect 3748 1060 3804 1062
rect 3828 1060 3884 1062
rect 3908 1060 3964 1062
rect 6550 1672 6606 1728
rect 6550 584 6606 640
rect 4328 570 4384 572
rect 4408 570 4464 572
rect 4488 570 4544 572
rect 4568 570 4624 572
rect 4328 518 4374 570
rect 4374 518 4384 570
rect 4408 518 4438 570
rect 4438 518 4450 570
rect 4450 518 4464 570
rect 4488 518 4502 570
rect 4502 518 4514 570
rect 4514 518 4544 570
rect 4568 518 4578 570
rect 4578 518 4624 570
rect 4328 516 4384 518
rect 4408 516 4464 518
rect 4488 516 4544 518
rect 4568 516 4624 518
<< metal3 >>
rect 7071 6808 7471 6928
rect 6269 6626 6335 6629
rect 7238 6626 7298 6808
rect 6269 6624 7298 6626
rect 6269 6568 6274 6624
rect 6330 6568 7298 6624
rect 6269 6566 7298 6568
rect 6269 6563 6335 6566
rect 3658 6560 3974 6561
rect 3658 6496 3664 6560
rect 3728 6496 3744 6560
rect 3808 6496 3824 6560
rect 3888 6496 3904 6560
rect 3968 6496 3974 6560
rect 3658 6495 3974 6496
rect 0 6082 400 6112
rect 4153 6082 4219 6085
rect 0 6080 4219 6082
rect 0 6024 4158 6080
rect 4214 6024 4219 6080
rect 0 6022 4219 6024
rect 0 5992 400 6022
rect 4153 6019 4219 6022
rect 6545 6082 6611 6085
rect 6545 6080 7298 6082
rect 6545 6024 6550 6080
rect 6606 6024 7298 6080
rect 6545 6022 7298 6024
rect 6545 6019 6611 6022
rect 4318 6016 4634 6017
rect 4318 5952 4324 6016
rect 4388 5952 4404 6016
rect 4468 5952 4484 6016
rect 4548 5952 4564 6016
rect 4628 5952 4634 6016
rect 4318 5951 4634 5952
rect 7238 5840 7298 6022
rect 7071 5720 7471 5840
rect 3658 5472 3974 5473
rect 3658 5408 3664 5472
rect 3728 5408 3744 5472
rect 3808 5408 3824 5472
rect 3888 5408 3904 5472
rect 3968 5408 3974 5472
rect 3658 5407 3974 5408
rect 6545 4994 6611 4997
rect 6545 4992 7298 4994
rect 6545 4936 6550 4992
rect 6606 4936 7298 4992
rect 6545 4934 7298 4936
rect 6545 4931 6611 4934
rect 4318 4928 4634 4929
rect 4318 4864 4324 4928
rect 4388 4864 4404 4928
rect 4468 4864 4484 4928
rect 4548 4864 4564 4928
rect 4628 4864 4634 4928
rect 4318 4863 4634 4864
rect 7238 4752 7298 4934
rect 7071 4632 7471 4752
rect 3658 4384 3974 4385
rect 3658 4320 3664 4384
rect 3728 4320 3744 4384
rect 3808 4320 3824 4384
rect 3888 4320 3904 4384
rect 3968 4320 3974 4384
rect 3658 4319 3974 4320
rect 6545 3906 6611 3909
rect 6545 3904 7298 3906
rect 6545 3848 6550 3904
rect 6606 3848 7298 3904
rect 6545 3846 7298 3848
rect 6545 3843 6611 3846
rect 4318 3840 4634 3841
rect 4318 3776 4324 3840
rect 4388 3776 4404 3840
rect 4468 3776 4484 3840
rect 4548 3776 4564 3840
rect 4628 3776 4634 3840
rect 4318 3775 4634 3776
rect 7238 3664 7298 3846
rect 0 3634 400 3664
rect 2773 3634 2839 3637
rect 0 3632 2839 3634
rect 0 3576 2778 3632
rect 2834 3576 2839 3632
rect 0 3574 2839 3576
rect 0 3544 400 3574
rect 2773 3571 2839 3574
rect 7071 3544 7471 3664
rect 3658 3296 3974 3297
rect 3658 3232 3664 3296
rect 3728 3232 3744 3296
rect 3808 3232 3824 3296
rect 3888 3232 3904 3296
rect 3968 3232 3974 3296
rect 3658 3231 3974 3232
rect 4318 2752 4634 2753
rect 4318 2688 4324 2752
rect 4388 2688 4404 2752
rect 4468 2688 4484 2752
rect 4548 2688 4564 2752
rect 4628 2688 4634 2752
rect 4318 2687 4634 2688
rect 6545 2546 6611 2549
rect 7071 2546 7471 2576
rect 6545 2544 7471 2546
rect 6545 2488 6550 2544
rect 6606 2488 7471 2544
rect 6545 2486 7471 2488
rect 6545 2483 6611 2486
rect 7054 2456 7471 2486
rect 7054 2452 7298 2456
rect 3658 2208 3974 2209
rect 3658 2144 3664 2208
rect 3728 2144 3744 2208
rect 3808 2144 3824 2208
rect 3888 2144 3904 2208
rect 3968 2144 3974 2208
rect 3658 2143 3974 2144
rect 6545 1730 6611 1733
rect 6545 1728 7298 1730
rect 6545 1672 6550 1728
rect 6606 1672 7298 1728
rect 6545 1670 7298 1672
rect 6545 1667 6611 1670
rect 4318 1664 4634 1665
rect 4318 1600 4324 1664
rect 4388 1600 4404 1664
rect 4468 1600 4484 1664
rect 4548 1600 4564 1664
rect 4628 1600 4634 1664
rect 4318 1599 4634 1600
rect 7238 1488 7298 1670
rect 7071 1368 7471 1488
rect 4797 1322 4863 1325
rect 2454 1320 4863 1322
rect 2454 1264 4802 1320
rect 4858 1264 4863 1320
rect 2454 1262 4863 1264
rect 0 1186 400 1216
rect 2454 1186 2514 1262
rect 4797 1259 4863 1262
rect 0 1126 2514 1186
rect 0 1096 400 1126
rect 3658 1120 3974 1121
rect 3658 1056 3664 1120
rect 3728 1056 3744 1120
rect 3808 1056 3824 1120
rect 3888 1056 3904 1120
rect 3968 1056 3974 1120
rect 3658 1055 3974 1056
rect 6545 642 6611 645
rect 6545 640 7298 642
rect 6545 584 6550 640
rect 6606 584 7298 640
rect 6545 582 7298 584
rect 6545 579 6611 582
rect 4318 576 4634 577
rect 4318 512 4324 576
rect 4388 512 4404 576
rect 4468 512 4484 576
rect 4548 512 4564 576
rect 4628 512 4634 576
rect 4318 511 4634 512
rect 7238 400 7298 582
rect 7071 280 7471 400
<< via3 >>
rect 3664 6556 3728 6560
rect 3664 6500 3668 6556
rect 3668 6500 3724 6556
rect 3724 6500 3728 6556
rect 3664 6496 3728 6500
rect 3744 6556 3808 6560
rect 3744 6500 3748 6556
rect 3748 6500 3804 6556
rect 3804 6500 3808 6556
rect 3744 6496 3808 6500
rect 3824 6556 3888 6560
rect 3824 6500 3828 6556
rect 3828 6500 3884 6556
rect 3884 6500 3888 6556
rect 3824 6496 3888 6500
rect 3904 6556 3968 6560
rect 3904 6500 3908 6556
rect 3908 6500 3964 6556
rect 3964 6500 3968 6556
rect 3904 6496 3968 6500
rect 4324 6012 4388 6016
rect 4324 5956 4328 6012
rect 4328 5956 4384 6012
rect 4384 5956 4388 6012
rect 4324 5952 4388 5956
rect 4404 6012 4468 6016
rect 4404 5956 4408 6012
rect 4408 5956 4464 6012
rect 4464 5956 4468 6012
rect 4404 5952 4468 5956
rect 4484 6012 4548 6016
rect 4484 5956 4488 6012
rect 4488 5956 4544 6012
rect 4544 5956 4548 6012
rect 4484 5952 4548 5956
rect 4564 6012 4628 6016
rect 4564 5956 4568 6012
rect 4568 5956 4624 6012
rect 4624 5956 4628 6012
rect 4564 5952 4628 5956
rect 3664 5468 3728 5472
rect 3664 5412 3668 5468
rect 3668 5412 3724 5468
rect 3724 5412 3728 5468
rect 3664 5408 3728 5412
rect 3744 5468 3808 5472
rect 3744 5412 3748 5468
rect 3748 5412 3804 5468
rect 3804 5412 3808 5468
rect 3744 5408 3808 5412
rect 3824 5468 3888 5472
rect 3824 5412 3828 5468
rect 3828 5412 3884 5468
rect 3884 5412 3888 5468
rect 3824 5408 3888 5412
rect 3904 5468 3968 5472
rect 3904 5412 3908 5468
rect 3908 5412 3964 5468
rect 3964 5412 3968 5468
rect 3904 5408 3968 5412
rect 4324 4924 4388 4928
rect 4324 4868 4328 4924
rect 4328 4868 4384 4924
rect 4384 4868 4388 4924
rect 4324 4864 4388 4868
rect 4404 4924 4468 4928
rect 4404 4868 4408 4924
rect 4408 4868 4464 4924
rect 4464 4868 4468 4924
rect 4404 4864 4468 4868
rect 4484 4924 4548 4928
rect 4484 4868 4488 4924
rect 4488 4868 4544 4924
rect 4544 4868 4548 4924
rect 4484 4864 4548 4868
rect 4564 4924 4628 4928
rect 4564 4868 4568 4924
rect 4568 4868 4624 4924
rect 4624 4868 4628 4924
rect 4564 4864 4628 4868
rect 3664 4380 3728 4384
rect 3664 4324 3668 4380
rect 3668 4324 3724 4380
rect 3724 4324 3728 4380
rect 3664 4320 3728 4324
rect 3744 4380 3808 4384
rect 3744 4324 3748 4380
rect 3748 4324 3804 4380
rect 3804 4324 3808 4380
rect 3744 4320 3808 4324
rect 3824 4380 3888 4384
rect 3824 4324 3828 4380
rect 3828 4324 3884 4380
rect 3884 4324 3888 4380
rect 3824 4320 3888 4324
rect 3904 4380 3968 4384
rect 3904 4324 3908 4380
rect 3908 4324 3964 4380
rect 3964 4324 3968 4380
rect 3904 4320 3968 4324
rect 4324 3836 4388 3840
rect 4324 3780 4328 3836
rect 4328 3780 4384 3836
rect 4384 3780 4388 3836
rect 4324 3776 4388 3780
rect 4404 3836 4468 3840
rect 4404 3780 4408 3836
rect 4408 3780 4464 3836
rect 4464 3780 4468 3836
rect 4404 3776 4468 3780
rect 4484 3836 4548 3840
rect 4484 3780 4488 3836
rect 4488 3780 4544 3836
rect 4544 3780 4548 3836
rect 4484 3776 4548 3780
rect 4564 3836 4628 3840
rect 4564 3780 4568 3836
rect 4568 3780 4624 3836
rect 4624 3780 4628 3836
rect 4564 3776 4628 3780
rect 3664 3292 3728 3296
rect 3664 3236 3668 3292
rect 3668 3236 3724 3292
rect 3724 3236 3728 3292
rect 3664 3232 3728 3236
rect 3744 3292 3808 3296
rect 3744 3236 3748 3292
rect 3748 3236 3804 3292
rect 3804 3236 3808 3292
rect 3744 3232 3808 3236
rect 3824 3292 3888 3296
rect 3824 3236 3828 3292
rect 3828 3236 3884 3292
rect 3884 3236 3888 3292
rect 3824 3232 3888 3236
rect 3904 3292 3968 3296
rect 3904 3236 3908 3292
rect 3908 3236 3964 3292
rect 3964 3236 3968 3292
rect 3904 3232 3968 3236
rect 4324 2748 4388 2752
rect 4324 2692 4328 2748
rect 4328 2692 4384 2748
rect 4384 2692 4388 2748
rect 4324 2688 4388 2692
rect 4404 2748 4468 2752
rect 4404 2692 4408 2748
rect 4408 2692 4464 2748
rect 4464 2692 4468 2748
rect 4404 2688 4468 2692
rect 4484 2748 4548 2752
rect 4484 2692 4488 2748
rect 4488 2692 4544 2748
rect 4544 2692 4548 2748
rect 4484 2688 4548 2692
rect 4564 2748 4628 2752
rect 4564 2692 4568 2748
rect 4568 2692 4624 2748
rect 4624 2692 4628 2748
rect 4564 2688 4628 2692
rect 3664 2204 3728 2208
rect 3664 2148 3668 2204
rect 3668 2148 3724 2204
rect 3724 2148 3728 2204
rect 3664 2144 3728 2148
rect 3744 2204 3808 2208
rect 3744 2148 3748 2204
rect 3748 2148 3804 2204
rect 3804 2148 3808 2204
rect 3744 2144 3808 2148
rect 3824 2204 3888 2208
rect 3824 2148 3828 2204
rect 3828 2148 3884 2204
rect 3884 2148 3888 2204
rect 3824 2144 3888 2148
rect 3904 2204 3968 2208
rect 3904 2148 3908 2204
rect 3908 2148 3964 2204
rect 3964 2148 3968 2204
rect 3904 2144 3968 2148
rect 4324 1660 4388 1664
rect 4324 1604 4328 1660
rect 4328 1604 4384 1660
rect 4384 1604 4388 1660
rect 4324 1600 4388 1604
rect 4404 1660 4468 1664
rect 4404 1604 4408 1660
rect 4408 1604 4464 1660
rect 4464 1604 4468 1660
rect 4404 1600 4468 1604
rect 4484 1660 4548 1664
rect 4484 1604 4488 1660
rect 4488 1604 4544 1660
rect 4544 1604 4548 1660
rect 4484 1600 4548 1604
rect 4564 1660 4628 1664
rect 4564 1604 4568 1660
rect 4568 1604 4624 1660
rect 4624 1604 4628 1660
rect 4564 1600 4628 1604
rect 3664 1116 3728 1120
rect 3664 1060 3668 1116
rect 3668 1060 3724 1116
rect 3724 1060 3728 1116
rect 3664 1056 3728 1060
rect 3744 1116 3808 1120
rect 3744 1060 3748 1116
rect 3748 1060 3804 1116
rect 3804 1060 3808 1116
rect 3744 1056 3808 1060
rect 3824 1116 3888 1120
rect 3824 1060 3828 1116
rect 3828 1060 3884 1116
rect 3884 1060 3888 1116
rect 3824 1056 3888 1060
rect 3904 1116 3968 1120
rect 3904 1060 3908 1116
rect 3908 1060 3964 1116
rect 3964 1060 3968 1116
rect 3904 1056 3968 1060
rect 4324 572 4388 576
rect 4324 516 4328 572
rect 4328 516 4384 572
rect 4384 516 4388 572
rect 4324 512 4388 516
rect 4404 572 4468 576
rect 4404 516 4408 572
rect 4408 516 4464 572
rect 4464 516 4468 572
rect 4404 512 4468 516
rect 4484 572 4548 576
rect 4484 516 4488 572
rect 4488 516 4544 572
rect 4544 516 4548 572
rect 4484 512 4548 516
rect 4564 572 4628 576
rect 4564 516 4568 572
rect 4568 516 4624 572
rect 4624 516 4628 572
rect 4564 512 4628 516
<< metal4 >>
rect 3656 6560 3976 6576
rect 3656 6496 3664 6560
rect 3728 6496 3744 6560
rect 3808 6496 3824 6560
rect 3888 6496 3904 6560
rect 3968 6496 3976 6560
rect 3656 5472 3976 6496
rect 3656 5408 3664 5472
rect 3728 5408 3744 5472
rect 3808 5408 3824 5472
rect 3888 5408 3904 5472
rect 3968 5408 3976 5472
rect 3656 4384 3976 5408
rect 3656 4320 3664 4384
rect 3728 4320 3744 4384
rect 3808 4320 3824 4384
rect 3888 4320 3904 4384
rect 3968 4320 3976 4384
rect 3656 3296 3976 4320
rect 3656 3232 3664 3296
rect 3728 3232 3744 3296
rect 3808 3232 3824 3296
rect 3888 3232 3904 3296
rect 3968 3232 3976 3296
rect 3656 2208 3976 3232
rect 3656 2144 3664 2208
rect 3728 2144 3744 2208
rect 3808 2144 3824 2208
rect 3888 2144 3904 2208
rect 3968 2144 3976 2208
rect 3656 1120 3976 2144
rect 3656 1056 3664 1120
rect 3728 1056 3744 1120
rect 3808 1056 3824 1120
rect 3888 1056 3904 1120
rect 3968 1056 3976 1120
rect 3656 496 3976 1056
rect 4316 6016 4636 6576
rect 4316 5952 4324 6016
rect 4388 5952 4404 6016
rect 4468 5952 4484 6016
rect 4548 5952 4564 6016
rect 4628 5952 4636 6016
rect 4316 4928 4636 5952
rect 4316 4864 4324 4928
rect 4388 4864 4404 4928
rect 4468 4864 4484 4928
rect 4548 4864 4564 4928
rect 4628 4864 4636 4928
rect 4316 3840 4636 4864
rect 4316 3776 4324 3840
rect 4388 3776 4404 3840
rect 4468 3776 4484 3840
rect 4548 3776 4564 3840
rect 4628 3776 4636 3840
rect 4316 2752 4636 3776
rect 4316 2688 4324 2752
rect 4388 2688 4404 2752
rect 4468 2688 4484 2752
rect 4548 2688 4564 2752
rect 4628 2688 4636 2752
rect 4316 1664 4636 2688
rect 4316 1600 4324 1664
rect 4388 1600 4404 1664
rect 4468 1600 4484 1664
rect 4548 1600 4564 1664
rect 4628 1600 4636 1664
rect 4316 576 4636 1600
rect 4316 512 4324 576
rect 4388 512 4404 576
rect 4468 512 4484 576
rect 4548 512 4564 576
rect 4628 512 4636 576
rect 4316 496 4636 512
use sky130_fd_sc_hd__and3_1  _09_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1755919380
transform 1 0 5244 0 -1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _10_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1755919380
transform -1 0 6532 0 -1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _11_
timestamp 1755919380
transform -1 0 5704 0 -1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _12_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1755919380
transform -1 0 5336 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__nor4_1  _13_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1755919380
transform -1 0 6348 0 -1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_4  _14_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1755919380
transform -1 0 6256 0 1 3808
box -38 -48 1326 592
use sky130_fd_sc_hd__a21o_2  _15_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1755919380
transform 1 0 4784 0 -1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _16_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1755919380
transform -1 0 6256 0 1 1632
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _17_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1755919380
transform -1 0 5796 0 1 1632
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _18_
timestamp 1755919380
transform 1 0 6348 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _19_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1755919380
transform 1 0 5796 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_4  _20_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1755919380
transform 1 0 4784 0 1 2720
box -38 -48 1602 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1755919380
transform 1 0 828 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15
timestamp 1755919380
transform 1 0 1932 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1755919380
transform 1 0 3036 0 1 544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29
timestamp 1755919380
transform 1 0 3220 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41
timestamp 1755919380
transform 1 0 4324 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1755919380
transform 1 0 5428 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1755919380
transform 1 0 5796 0 1 544
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3
timestamp 1755919380
transform 1 0 828 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_15
timestamp 1755919380
transform 1 0 1932 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_27
timestamp 1755919380
transform 1 0 3036 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_39
timestamp 1755919380
transform 1 0 4140 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1755919380
transform 1 0 5244 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1755919380
transform 1 0 5612 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_57 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1755919380
transform 1 0 5796 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_65
timestamp 1755919380
transform 1 0 6532 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 1755919380
transform 1 0 828 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1755919380
transform 1 0 1932 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1755919380
transform 1 0 3036 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1755919380
transform 1 0 3220 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_41
timestamp 1755919380
transform 1 0 4324 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_62
timestamp 1755919380
transform 1 0 6256 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1755919380
transform 1 0 828 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1755919380
transform 1 0 1932 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1755919380
transform 1 0 3036 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 1755919380
transform 1 0 4140 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_57
timestamp 1755919380
transform 1 0 5796 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1755919380
transform 1 0 828 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1755919380
transform 1 0 1932 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1755919380
transform 1 0 3036 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1755919380
transform 1 0 3220 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_41
timestamp 1755919380
transform 1 0 4324 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_45
timestamp 1755919380
transform 1 0 4692 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1755919380
transform 1 0 828 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1755919380
transform 1 0 1932 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_27
timestamp 1755919380
transform 1 0 3036 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_39
timestamp 1755919380
transform 1 0 4140 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_45
timestamp 1755919380
transform 1 0 4692 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_5_53
timestamp 1755919380
transform 1 0 5428 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_57
timestamp 1755919380
transform 1 0 5796 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_65
timestamp 1755919380
transform 1 0 6532 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1755919380
transform 1 0 828 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1755919380
transform 1 0 1932 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1755919380
transform 1 0 3036 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1755919380
transform 1 0 3220 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_41
timestamp 1755919380
transform 1 0 4324 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_47
timestamp 1755919380
transform 1 0 4876 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_62
timestamp 1755919380
transform 1 0 6256 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1755919380
transform 1 0 828 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1755919380
transform 1 0 1932 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1755919380
transform 1 0 3036 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_39
timestamp 1755919380
transform 1 0 4140 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1755919380
transform 1 0 828 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1755919380
transform 1 0 1932 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1755919380
transform 1 0 3036 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1755919380
transform 1 0 3220 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1755919380
transform 1 0 4324 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_53
timestamp 1755919380
transform 1 0 5428 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_61 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1755919380
transform 1 0 6164 0 1 4896
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1755919380
transform 1 0 828 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_15
timestamp 1755919380
transform 1 0 1932 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_27
timestamp 1755919380
transform 1 0 3036 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_39
timestamp 1755919380
transform 1 0 4140 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp 1755919380
transform 1 0 5244 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1755919380
transform 1 0 5612 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_57
timestamp 1755919380
transform 1 0 5796 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_65
timestamp 1755919380
transform 1 0 6532 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1755919380
transform 1 0 828 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1755919380
transform 1 0 1932 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1755919380
transform 1 0 3036 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1755919380
transform 1 0 3220 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1755919380
transform 1 0 4324 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_10_53
timestamp 1755919380
transform 1 0 5428 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_57
timestamp 1755919380
transform 1 0 5796 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input1 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1755919380
transform -1 0 6348 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input2
timestamp 1755919380
transform -1 0 6624 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1755919380
transform 1 0 6348 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1755919380
transform 1 0 6348 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input5
timestamp 1755919380
transform -1 0 6624 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input6
timestamp 1755919380
transform -1 0 6624 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input7
timestamp 1755919380
transform -1 0 6624 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  max_cap8
timestamp 1755919380
transform 1 0 6348 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_11
timestamp 1755919380
transform 1 0 552 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 1755919380
transform -1 0 6900 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_12
timestamp 1755919380
transform 1 0 552 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 1755919380
transform -1 0 6900 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_13
timestamp 1755919380
transform 1 0 552 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 1755919380
transform -1 0 6900 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_14
timestamp 1755919380
transform 1 0 552 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 1755919380
transform -1 0 6900 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_15
timestamp 1755919380
transform 1 0 552 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 1755919380
transform -1 0 6900 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_16
timestamp 1755919380
transform 1 0 552 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 1755919380
transform -1 0 6900 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_17
timestamp 1755919380
transform 1 0 552 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 1755919380
transform -1 0 6900 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_18
timestamp 1755919380
transform 1 0 552 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 1755919380
transform -1 0 6900 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_19
timestamp 1755919380
transform 1 0 552 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 1755919380
transform -1 0 6900 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_20
timestamp 1755919380
transform 1 0 552 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 1755919380
transform -1 0 6900 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_21
timestamp 1755919380
transform 1 0 552 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 1755919380
transform -1 0 6900 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_22 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1755919380
transform 1 0 3128 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_23
timestamp 1755919380
transform 1 0 5704 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_24
timestamp 1755919380
transform 1 0 5704 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_25
timestamp 1755919380
transform 1 0 3128 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_26
timestamp 1755919380
transform 1 0 5704 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_27
timestamp 1755919380
transform 1 0 3128 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_28
timestamp 1755919380
transform 1 0 5704 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_29
timestamp 1755919380
transform 1 0 3128 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_30
timestamp 1755919380
transform 1 0 5704 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_31
timestamp 1755919380
transform 1 0 3128 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_32
timestamp 1755919380
transform 1 0 5704 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_33
timestamp 1755919380
transform 1 0 3128 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_34
timestamp 1755919380
transform 1 0 5704 0 1 5984
box -38 -48 130 592
<< labels >>
flabel metal4 s 4316 496 4636 6576 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 3656 496 3976 6576 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal2 s 3698 0 3754 400 0 FreeSans 224 90 0 0 clk
port 2 nsew signal input
flabel metal3 s 0 1096 400 1216 0 FreeSans 480 0 0 0 o0
port 3 nsew signal output
flabel metal3 s 0 3544 400 3664 0 FreeSans 480 0 0 0 o1
port 4 nsew signal output
flabel metal3 s 0 5992 400 6112 0 FreeSans 480 0 0 0 o2
port 5 nsew signal output
flabel metal3 s 7071 6808 7471 6928 0 FreeSans 480 0 0 0 t0
port 6 nsew signal input
flabel metal3 s 7071 5720 7471 5840 0 FreeSans 480 0 0 0 t1
port 7 nsew signal input
flabel metal3 s 7071 4632 7471 4752 0 FreeSans 480 0 0 0 t2
port 8 nsew signal input
flabel metal3 s 7071 3544 7471 3664 0 FreeSans 480 0 0 0 t3
port 9 nsew signal input
flabel metal3 s 7071 2456 7471 2576 0 FreeSans 480 0 0 0 t4
port 10 nsew signal input
flabel metal3 s 7071 1368 7471 1488 0 FreeSans 480 0 0 0 t5
port 11 nsew signal input
flabel metal3 s 7071 280 7471 400 0 FreeSans 480 0 0 0 t6
port 12 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 7471 7455
<< end >>
