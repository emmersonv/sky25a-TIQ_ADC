** sch_path: /foss/designs/analog-circuit-design/sky25a-TIQ_ADC/xschem/INVERTER_SIZES/inverter_p3_n3o5_symsch.sch
.subckt inverter_p3_n3o5_symsch Vout Vin VDPWR VGND
*.PININFO Vout:O Vin:I VDPWR:B VGND:B
x1 VDPWR Vout Vin VGND inverter_p3_n3o5
.ends

* expanding   symbol:  /foss/designs/analog-circuit-design/sky25a-TIQ_ADC/xschem/INVERTER_SIZES/inverter_p3_n3o5.sym # of pins=4
** sym_path: /foss/designs/analog-circuit-design/sky25a-TIQ_ADC/xschem/INVERTER_SIZES/inverter_p3_n3o5.sym
** sch_path: /foss/designs/analog-circuit-design/sky25a-TIQ_ADC/xschem/INVERTER_SIZES/inverter_p3_n3o5.sch
.subckt inverter_p3_n3o5 VDPWR Vout Vin VGND
*.PININFO Vout:O Vin:I VDPWR:B VGND:B
XM1 Vout Vin VGND VGND sky130_fd_pr__nfet_01v8 L=0.15 W=3.5 nf=1 m=1
XM2 Vout Vin VDPWR VDPWR sky130_fd_pr__pfet_01v8 L=0.15 W=3 nf=1 m=1
.ends

