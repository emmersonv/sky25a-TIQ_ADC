magic
tech sky130A
magscale 1 2
timestamp 1756008383
<< nwell >>
rect -80 656 334 2996
<< pwell >>
rect -108 -1026 360 -774
<< psubdiff >>
rect -82 -833 334 -800
rect -82 -867 -3 -833
rect 31 -867 89 -833
rect 123 -867 181 -833
rect 215 -867 273 -833
rect 307 -867 334 -833
rect -82 -925 334 -867
rect -82 -959 -3 -925
rect 31 -959 89 -925
rect 123 -959 181 -925
rect 215 -959 273 -925
rect 307 -959 334 -925
rect -82 -1000 334 -959
<< nsubdiff >>
rect 0 2929 252 2960
rect 0 2895 31 2929
rect 65 2895 123 2929
rect 157 2895 252 2929
rect 0 2837 252 2895
rect 0 2803 31 2837
rect 65 2803 123 2837
rect 157 2803 252 2837
rect 0 2760 252 2803
<< psubdiffcont >>
rect -3 -867 31 -833
rect 89 -867 123 -833
rect 181 -867 215 -833
rect 273 -867 307 -833
rect -3 -959 31 -925
rect 89 -959 123 -925
rect 181 -959 215 -925
rect 273 -959 307 -925
<< nsubdiffcont >>
rect 31 2895 65 2929
rect 123 2895 157 2929
rect 31 2803 65 2837
rect 123 2803 157 2837
<< poly >>
rect -80 676 -14 692
rect -80 642 -64 676
rect -30 656 -14 676
rect 62 656 188 662
rect -30 644 188 656
rect -30 642 62 644
rect -80 626 62 642
<< polycont >>
rect -64 642 -30 676
<< locali >>
rect -80 2929 334 2946
rect -80 2895 -61 2929
rect -27 2895 31 2929
rect 65 2895 123 2929
rect 157 2895 215 2929
rect 249 2895 334 2929
rect -80 2837 334 2895
rect -80 2803 -61 2837
rect -27 2803 31 2837
rect 65 2803 123 2837
rect 157 2803 215 2837
rect 249 2803 334 2837
rect -80 2774 334 2803
rect 12 2222 46 2774
rect 204 2222 238 2774
rect -80 676 -14 692
rect -80 642 -64 676
rect -30 642 -14 676
rect -80 626 -14 642
rect 108 666 142 714
rect 268 676 334 692
rect 268 666 284 676
rect 108 642 284 666
rect 318 642 334 676
rect 108 626 334 642
rect 108 592 142 626
rect 12 -816 46 84
rect 204 -816 238 84
rect -80 -833 334 -816
rect -80 -867 -3 -833
rect 31 -867 89 -833
rect 123 -867 181 -833
rect 215 -867 273 -833
rect 307 -867 334 -833
rect -80 -925 334 -867
rect -80 -959 -3 -925
rect 31 -959 89 -925
rect 123 -959 181 -925
rect 215 -959 273 -925
rect 307 -959 334 -925
rect -80 -984 334 -959
<< viali >>
rect -61 2895 -27 2929
rect 31 2895 65 2929
rect 123 2895 157 2929
rect 215 2895 249 2929
rect -61 2803 -27 2837
rect 31 2803 65 2837
rect 123 2803 157 2837
rect 215 2803 249 2837
rect -64 642 -30 676
rect 284 642 318 676
rect -3 -867 31 -833
rect 89 -867 123 -833
rect 181 -867 215 -833
rect 273 -867 307 -833
rect -3 -959 31 -925
rect 89 -959 123 -925
rect 181 -959 215 -925
rect 273 -959 307 -925
<< metal1 >>
rect -80 2929 334 2946
rect -80 2895 -61 2929
rect -27 2895 31 2929
rect 65 2895 123 2929
rect 157 2895 215 2929
rect 249 2895 334 2929
rect -80 2837 334 2895
rect -80 2803 -61 2837
rect -27 2803 31 2837
rect 65 2803 123 2837
rect 157 2803 215 2837
rect 249 2803 334 2837
rect -80 2774 334 2803
rect -80 676 -14 692
rect -80 642 -64 676
rect -30 642 -14 676
rect -80 626 -14 642
rect 268 676 334 692
rect 268 642 284 676
rect 318 642 334 676
rect 268 626 334 642
rect -80 -833 334 -816
rect -80 -867 -3 -833
rect 31 -867 89 -833
rect 123 -867 181 -833
rect 215 -867 273 -833
rect 307 -867 334 -833
rect -80 -925 334 -867
rect -80 -959 -3 -925
rect 31 -959 89 -925
rect 123 -959 181 -925
rect 215 -959 273 -925
rect 307 -959 334 -925
rect -80 -984 334 -959
use sky130_fd_pr__nfet_01v8_V2VUT3  sky130_fd_pr__nfet_01v8_V2VUT3_0
timestamp 1756008383
transform 1 0 125 0 1 338
box -151 -276 151 306
use sky130_fd_pr__pfet_01v8_7QKTNL  sky130_fd_pr__pfet_01v8_7QKTNL_0
timestamp 1756008383
transform 1 0 125 0 1 1468
box -161 -812 161 812
<< end >>
