magic
tech sky130A
magscale 1 2
timestamp 1755919380
<< error_s >>
rect -248 318 -232 470
rect -196 318 22 572
rect 212 318 430 572
rect -248 302 22 318
rect -196 294 -92 302
rect 326 294 430 318
rect 466 318 482 470
rect 466 302 634 318
<< nwell >>
rect -196 2418 430 2646
rect -148 2410 -114 2418
rect 44 2410 78 2418
rect 156 2410 190 2418
rect 348 2410 382 2418
rect -196 2394 430 2410
rect -148 2360 -114 2394
rect 44 2360 78 2394
rect 156 2360 190 2394
rect 348 2360 382 2394
rect -248 302 -232 318
rect 28 300 206 330
rect 466 302 482 318
<< psubdiff >>
rect -248 -1182 470 -1150
rect -248 -1218 -236 -1182
rect -200 -1218 -144 -1182
rect -108 -1218 -52 -1182
rect -16 -1218 40 -1182
rect 76 -1218 132 -1182
rect 168 -1218 224 -1182
rect 260 -1218 316 -1182
rect 352 -1218 408 -1182
rect 444 -1218 470 -1182
rect -248 -1274 470 -1218
rect -248 -1310 -236 -1274
rect -200 -1310 -144 -1274
rect -108 -1310 -52 -1274
rect -16 -1310 40 -1274
rect 76 -1310 132 -1274
rect 168 -1310 224 -1274
rect 260 -1310 316 -1274
rect 352 -1310 408 -1274
rect 444 -1310 470 -1274
rect -248 -1350 470 -1310
<< nsubdiff >>
rect -160 2580 394 2610
rect -160 2544 -110 2580
rect -74 2544 -18 2580
rect 18 2544 74 2580
rect 110 2544 166 2580
rect 202 2544 258 2580
rect 294 2544 350 2580
rect 386 2544 394 2580
rect -160 2488 394 2544
rect -160 2452 -110 2488
rect -74 2452 -18 2488
rect 18 2452 74 2488
rect 110 2452 166 2488
rect 202 2452 258 2488
rect 294 2452 350 2488
rect 386 2452 394 2488
rect -160 2410 394 2452
<< psubdiffcont >>
rect -236 -1218 -200 -1182
rect -144 -1218 -108 -1182
rect -52 -1218 -16 -1182
rect 40 -1218 76 -1182
rect 132 -1218 168 -1182
rect 224 -1218 260 -1182
rect 316 -1218 352 -1182
rect 408 -1218 444 -1182
rect -236 -1310 -200 -1274
rect -144 -1310 -108 -1274
rect -52 -1310 -16 -1274
rect 40 -1310 76 -1274
rect 132 -1310 168 -1274
rect 224 -1310 260 -1274
rect 316 -1310 352 -1274
rect 408 -1310 444 -1274
<< nsubdiffcont >>
rect -110 2544 -74 2580
rect -18 2544 18 2580
rect 74 2544 110 2580
rect 166 2544 202 2580
rect 258 2544 294 2580
rect 350 2544 386 2580
rect -110 2452 -74 2488
rect -18 2452 18 2488
rect 74 2452 110 2488
rect 166 2452 202 2488
rect 258 2452 294 2488
rect 350 2452 386 2488
<< poly >>
rect -248 326 -182 342
rect -248 292 -232 326
rect -198 306 -182 326
rect 28 306 206 330
rect -198 300 206 306
rect -198 292 332 300
rect -248 276 332 292
rect 58 252 88 276
<< polycont >>
rect -232 292 -198 326
<< locali >>
rect -248 2580 516 2596
rect -248 2544 -202 2580
rect -166 2544 -110 2580
rect -74 2544 -18 2580
rect 18 2544 74 2580
rect 110 2544 166 2580
rect 202 2544 258 2580
rect 294 2544 350 2580
rect 386 2544 516 2580
rect -248 2488 516 2544
rect -248 2452 -202 2488
rect -166 2452 -110 2488
rect -74 2452 -18 2488
rect 18 2452 74 2488
rect 110 2452 166 2488
rect 202 2452 258 2488
rect 294 2452 350 2488
rect 386 2452 516 2488
rect -248 2424 516 2452
rect -148 2360 -114 2424
rect 44 2360 78 2424
rect 156 2360 190 2424
rect 348 2360 382 2424
rect -248 326 -182 342
rect -248 292 -232 326
rect -198 292 -182 326
rect -248 276 -182 292
rect -52 316 -18 368
rect 252 316 286 352
rect 416 326 482 342
rect 416 316 432 326
rect -52 292 432 316
rect 466 292 482 326
rect -52 276 482 292
rect 100 230 134 276
rect 12 -1166 46 22
rect -248 -1182 470 -1166
rect -248 -1218 -236 -1182
rect -200 -1218 -144 -1182
rect -108 -1218 -52 -1182
rect -16 -1218 40 -1182
rect 76 -1218 132 -1182
rect 168 -1218 224 -1182
rect 260 -1218 316 -1182
rect 352 -1218 408 -1182
rect 444 -1218 470 -1182
rect -248 -1274 470 -1218
rect -248 -1310 -236 -1274
rect -200 -1310 -144 -1274
rect -108 -1310 -52 -1274
rect -16 -1310 40 -1274
rect 76 -1310 132 -1274
rect 168 -1310 224 -1274
rect 260 -1310 316 -1274
rect 352 -1310 408 -1274
rect 444 -1310 470 -1274
rect -248 -1334 470 -1310
<< viali >>
rect -202 2544 -166 2580
rect -110 2544 -74 2580
rect -18 2544 18 2580
rect 74 2544 110 2580
rect 166 2544 202 2580
rect 258 2544 294 2580
rect 350 2544 386 2580
rect -202 2452 -166 2488
rect -110 2452 -74 2488
rect -18 2452 18 2488
rect 74 2452 110 2488
rect 166 2452 202 2488
rect 258 2452 294 2488
rect 350 2452 386 2488
rect -232 292 -198 326
rect 432 292 466 326
rect -236 -1218 -200 -1182
rect -144 -1218 -108 -1182
rect -52 -1218 -16 -1182
rect 40 -1218 76 -1182
rect 132 -1218 168 -1182
rect 224 -1218 260 -1182
rect 316 -1218 352 -1182
rect 408 -1218 444 -1182
rect -236 -1310 -200 -1274
rect -144 -1310 -108 -1274
rect -52 -1310 -16 -1274
rect 40 -1310 76 -1274
rect 132 -1310 168 -1274
rect 224 -1310 260 -1274
rect 316 -1310 352 -1274
rect 408 -1310 444 -1274
<< metal1 >>
rect -248 2580 516 2596
rect -248 2544 -202 2580
rect -166 2544 -110 2580
rect -74 2544 -18 2580
rect 18 2544 74 2580
rect 110 2544 166 2580
rect 202 2544 258 2580
rect 294 2544 350 2580
rect 386 2544 516 2580
rect -248 2488 516 2544
rect -248 2452 -202 2488
rect -166 2452 -110 2488
rect -74 2452 -18 2488
rect 18 2452 74 2488
rect 110 2452 166 2488
rect 202 2452 258 2488
rect 294 2452 350 2488
rect 386 2452 516 2488
rect -248 2424 516 2452
rect -248 326 -182 342
rect -248 292 -232 326
rect -198 292 -182 326
rect -248 276 -182 292
rect 416 326 482 342
rect 416 292 432 326
rect 466 292 482 326
rect 416 276 482 292
rect -248 -1182 470 -1166
rect -248 -1218 -236 -1182
rect -200 -1218 -144 -1182
rect -108 -1218 -52 -1182
rect -16 -1218 40 -1182
rect 76 -1218 132 -1182
rect 168 -1218 224 -1182
rect 260 -1218 316 -1182
rect 352 -1218 408 -1182
rect 444 -1218 470 -1182
rect -248 -1274 470 -1218
rect -248 -1310 -236 -1274
rect -200 -1310 -144 -1274
rect -108 -1310 -52 -1274
rect -16 -1310 40 -1274
rect 76 -1310 132 -1274
rect 168 -1310 224 -1274
rect 260 -1310 316 -1274
rect 352 -1310 408 -1274
rect 444 -1310 470 -1274
rect -248 -1334 470 -1310
use sky130_fd_pr__nfet_01v8_QDUU3W  sky130_fd_pr__nfet_01v8_QDUU3W_0
timestamp 1755919380
transform 1 0 73 0 1 126
box -73 -126 73 126
use sky130_fd_pr__pfet_01v8_WELYR5  sky130_fd_pr__pfet_01v8_WELYR5_0
timestamp 1755919380
transform 1 0 -35 0 1 1356
box -161 -1062 161 1062
use sky130_fd_pr__pfet_01v8_WELYR5  sky130_fd_pr__pfet_01v8_WELYR5_1
timestamp 1755919380
transform 1 0 269 0 1 1356
box -161 -1062 161 1062
<< end >>
