magic
tech sky130A
magscale 1 2
timestamp 1756008383
<< error_s >>
rect 4640 4300 4840 4458
rect 4876 4300 5008 4468
rect 4640 4264 5008 4300
rect 4840 4240 5008 4264
rect 4640 4204 5008 4240
rect 4640 4168 4840 4204
<< poly >>
rect 740 6321 774 6322
rect 740 6286 774 6287
rect 740 5337 774 5338
rect 740 5302 774 5303
rect 740 4351 774 4352
rect 740 4316 774 4317
rect 740 3367 774 3368
rect 740 3332 774 3333
rect 740 2383 774 2384
rect 740 2348 774 2349
rect 740 1399 774 1400
rect 740 1364 774 1365
rect 740 415 774 416
rect 740 380 774 381
<< polycont >>
rect 740 6287 774 6321
rect 740 5303 774 5337
rect 740 4317 774 4351
rect 740 3333 774 3367
rect 740 2349 774 2383
rect 740 1365 774 1399
rect 740 381 774 415
<< locali >>
rect 4 6282 52 6322
rect 724 6321 790 6338
rect 724 6287 740 6321
rect 774 6287 790 6321
rect 724 6270 790 6287
rect 896 5815 1064 5882
rect 896 5781 921 5815
rect 955 5781 1064 5815
rect 4 5298 52 5338
rect 724 5337 790 5354
rect 724 5303 740 5337
rect 774 5303 790 5337
rect 724 5286 790 5303
rect 4 4312 52 4352
rect 724 4351 790 4368
rect 724 4317 740 4351
rect 774 4317 790 4351
rect 724 4300 790 4317
rect 4 3328 52 3368
rect 724 3367 790 3384
rect 724 3333 740 3367
rect 774 3333 790 3367
rect 724 3316 790 3333
rect 4 2344 52 2384
rect 724 2383 790 2400
rect 724 2349 740 2383
rect 774 2349 790 2383
rect 724 2332 790 2349
rect 4 1360 52 1400
rect 724 1399 790 1416
rect 724 1365 740 1399
rect 774 1365 790 1399
rect 724 1348 790 1365
rect 896 758 1064 5781
rect 4654 1787 4826 5882
rect 4654 1753 4775 1787
rect 4809 1753 4826 1787
rect 4654 760 4826 1753
rect 4 376 52 416
rect 724 415 790 432
rect 724 381 740 415
rect 774 381 790 415
rect 724 364 790 381
<< viali >>
rect 740 6287 774 6321
rect 921 5781 955 5815
rect 740 5303 774 5337
rect 740 4317 774 4351
rect 740 3333 774 3367
rect 740 2349 774 2383
rect 740 1365 774 1399
rect 4775 1753 4809 1787
rect 740 381 774 415
<< metal1 >>
rect -260 6642 4 6814
rect 790 6642 4826 6818
rect -260 5832 -110 6642
rect 724 6331 790 6338
rect 724 6279 731 6331
rect 783 6279 790 6331
rect 724 6270 790 6279
rect 790 5924 1082 6092
rect 880 5882 1082 5924
rect -260 5660 4 5832
rect 896 5815 1064 5882
rect 896 5781 921 5815
rect 955 5781 1064 5815
rect -260 4844 -110 5660
rect 724 5347 790 5354
rect 724 5295 731 5347
rect 783 5295 790 5347
rect 724 5286 790 5295
rect 896 5106 1064 5781
rect 790 4938 1064 5106
rect -260 4672 4 4844
rect -260 3860 -110 4672
rect 724 4359 790 4368
rect 724 4307 731 4359
rect 783 4307 790 4359
rect 724 4300 790 4307
rect 896 4122 1064 4938
rect 792 3954 1064 4122
rect -260 3688 6 3860
rect -260 2876 -110 3688
rect 724 3377 790 3384
rect 724 3325 731 3377
rect 783 3325 790 3377
rect 724 3316 790 3325
rect 896 3136 1064 3954
rect 790 2968 1064 3136
rect -260 2704 4 2876
rect -260 1892 -110 2704
rect 724 2393 790 2400
rect 724 2341 731 2393
rect 783 2341 790 2393
rect 724 2332 790 2341
rect 896 2154 1064 2968
rect 790 1986 1064 2154
rect -260 1720 4 1892
rect -260 908 -110 1720
rect 724 1409 790 1416
rect 724 1357 731 1409
rect 783 1357 790 1409
rect 724 1348 790 1357
rect 896 1170 1064 1986
rect 790 1002 1064 1170
rect -260 736 2 908
rect 724 425 790 432
rect 724 373 731 425
rect 783 373 790 425
rect 724 364 790 373
rect 896 184 1064 1002
rect 4654 1787 4826 6642
rect 4654 1753 4775 1787
rect 4809 1753 4826 1787
rect 4654 760 4826 1753
rect 790 16 1064 184
<< via1 >>
rect 731 6321 783 6331
rect 731 6287 740 6321
rect 740 6287 774 6321
rect 774 6287 783 6321
rect 731 6279 783 6287
rect 731 5337 783 5347
rect 731 5303 740 5337
rect 740 5303 774 5337
rect 774 5303 783 5337
rect 731 5295 783 5303
rect 731 4351 783 4359
rect 731 4317 740 4351
rect 740 4317 774 4351
rect 774 4317 783 4351
rect 731 4307 783 4317
rect 731 3367 783 3377
rect 731 3333 740 3367
rect 740 3333 774 3367
rect 774 3333 783 3367
rect 731 3325 783 3333
rect 731 2383 783 2393
rect 731 2349 740 2383
rect 740 2349 774 2383
rect 774 2349 783 2383
rect 731 2341 783 2349
rect 731 1399 783 1409
rect 731 1365 740 1399
rect 740 1365 774 1399
rect 774 1365 783 1399
rect 731 1357 783 1365
rect 731 415 783 425
rect 731 381 740 415
rect 740 381 774 415
rect 774 381 783 415
rect 731 373 783 381
<< metal2 >>
rect 724 6331 2464 6338
rect 724 6279 731 6331
rect 783 6279 2464 6331
rect 724 6270 2464 6279
rect 724 5347 2370 5354
rect 724 5295 731 5347
rect 783 5295 2370 5347
rect 724 5286 2370 5295
rect 2304 4446 2370 5286
rect 2398 5054 2464 6270
rect 2398 4988 2572 5054
rect 2304 4380 2572 4446
rect 724 4359 2276 4368
rect 724 4307 731 4359
rect 783 4307 2276 4359
rect 724 4300 2276 4307
rect 2210 3838 2276 4300
rect 2210 3772 2572 3838
rect 724 3377 2572 3390
rect 724 3325 731 3377
rect 783 3325 2572 3377
rect 724 3324 2572 3325
rect 724 3316 790 3324
rect 2398 2880 2506 2946
rect 2398 2400 2464 2880
rect 724 2393 2464 2400
rect 724 2341 731 2393
rect 783 2341 2464 2393
rect 724 2332 2464 2341
rect 2398 2116 2506 2182
rect 2398 1416 2464 2116
rect 2602 2032 2636 5830
rect 724 1409 2464 1416
rect 724 1357 731 1409
rect 783 1357 2464 1409
rect 724 1348 2464 1357
rect 2508 432 2574 760
rect 724 425 2574 432
rect 724 373 731 425
rect 783 373 2574 425
rect 724 364 2574 373
use gain_stage_7  gain_stage_7_0
timestamp 1756008383
transform -1 0 790 0 1 5906
box -28 -5932 814 958
use tiq_adc_7  tiq_adc_7_0
timestamp 1756008383
transform 1 0 880 0 1 760
box -26 -26 4128 5148
<< labels >>
rlabel metal1 s 2368 6642 2532 6818 4 VDPWR
port 1 nsew
rlabel metal1 s 896 16 1058 172 4 VGND
port 2 nsew
rlabel metal2 s 2602 3558 2636 3604 4 Vin
port 3 nsew
rlabel locali s 10 6290 36 6314 4 t0
port 4 nsew
rlabel locali s 12 5306 38 5330 4 t1
port 5 nsew
rlabel locali s 10 4318 36 4342 4 t2
port 6 nsew
rlabel locali s 10 3336 36 3360 4 t3
port 7 nsew
rlabel locali s 10 2352 36 2376 4 t4
port 8 nsew
rlabel locali s 10 1368 36 1392 4 t5
port 9 nsew
rlabel locali s 8 384 34 408 4 t6
port 10 nsew
<< end >>
