magic
tech sky130A
magscale 1 2
timestamp 1756008383
<< nwell >>
rect -161 -1062 161 1062
<< pmos >>
rect -63 -1000 -33 1000
rect 33 -1000 63 1000
<< pdiff >>
rect -125 969 -63 1000
rect -125 935 -113 969
rect -79 935 -63 969
rect -125 901 -63 935
rect -125 867 -113 901
rect -79 867 -63 901
rect -125 833 -63 867
rect -125 799 -113 833
rect -79 799 -63 833
rect -125 765 -63 799
rect -125 731 -113 765
rect -79 731 -63 765
rect -125 697 -63 731
rect -125 663 -113 697
rect -79 663 -63 697
rect -125 629 -63 663
rect -125 595 -113 629
rect -79 595 -63 629
rect -125 561 -63 595
rect -125 527 -113 561
rect -79 527 -63 561
rect -125 493 -63 527
rect -125 459 -113 493
rect -79 459 -63 493
rect -125 425 -63 459
rect -125 391 -113 425
rect -79 391 -63 425
rect -125 357 -63 391
rect -125 323 -113 357
rect -79 323 -63 357
rect -125 289 -63 323
rect -125 255 -113 289
rect -79 255 -63 289
rect -125 221 -63 255
rect -125 187 -113 221
rect -79 187 -63 221
rect -125 153 -63 187
rect -125 119 -113 153
rect -79 119 -63 153
rect -125 85 -63 119
rect -125 51 -113 85
rect -79 51 -63 85
rect -125 17 -63 51
rect -125 -17 -113 17
rect -79 -17 -63 17
rect -125 -51 -63 -17
rect -125 -85 -113 -51
rect -79 -85 -63 -51
rect -125 -119 -63 -85
rect -125 -153 -113 -119
rect -79 -153 -63 -119
rect -125 -187 -63 -153
rect -125 -221 -113 -187
rect -79 -221 -63 -187
rect -125 -255 -63 -221
rect -125 -289 -113 -255
rect -79 -289 -63 -255
rect -125 -323 -63 -289
rect -125 -357 -113 -323
rect -79 -357 -63 -323
rect -125 -391 -63 -357
rect -125 -425 -113 -391
rect -79 -425 -63 -391
rect -125 -459 -63 -425
rect -125 -493 -113 -459
rect -79 -493 -63 -459
rect -125 -527 -63 -493
rect -125 -561 -113 -527
rect -79 -561 -63 -527
rect -125 -595 -63 -561
rect -125 -629 -113 -595
rect -79 -629 -63 -595
rect -125 -663 -63 -629
rect -125 -697 -113 -663
rect -79 -697 -63 -663
rect -125 -731 -63 -697
rect -125 -765 -113 -731
rect -79 -765 -63 -731
rect -125 -799 -63 -765
rect -125 -833 -113 -799
rect -79 -833 -63 -799
rect -125 -867 -63 -833
rect -125 -901 -113 -867
rect -79 -901 -63 -867
rect -125 -935 -63 -901
rect -125 -969 -113 -935
rect -79 -969 -63 -935
rect -125 -1000 -63 -969
rect -33 969 33 1000
rect -33 935 -17 969
rect 17 935 33 969
rect -33 901 33 935
rect -33 867 -17 901
rect 17 867 33 901
rect -33 833 33 867
rect -33 799 -17 833
rect 17 799 33 833
rect -33 765 33 799
rect -33 731 -17 765
rect 17 731 33 765
rect -33 697 33 731
rect -33 663 -17 697
rect 17 663 33 697
rect -33 629 33 663
rect -33 595 -17 629
rect 17 595 33 629
rect -33 561 33 595
rect -33 527 -17 561
rect 17 527 33 561
rect -33 493 33 527
rect -33 459 -17 493
rect 17 459 33 493
rect -33 425 33 459
rect -33 391 -17 425
rect 17 391 33 425
rect -33 357 33 391
rect -33 323 -17 357
rect 17 323 33 357
rect -33 289 33 323
rect -33 255 -17 289
rect 17 255 33 289
rect -33 221 33 255
rect -33 187 -17 221
rect 17 187 33 221
rect -33 153 33 187
rect -33 119 -17 153
rect 17 119 33 153
rect -33 85 33 119
rect -33 51 -17 85
rect 17 51 33 85
rect -33 17 33 51
rect -33 -17 -17 17
rect 17 -17 33 17
rect -33 -51 33 -17
rect -33 -85 -17 -51
rect 17 -85 33 -51
rect -33 -119 33 -85
rect -33 -153 -17 -119
rect 17 -153 33 -119
rect -33 -187 33 -153
rect -33 -221 -17 -187
rect 17 -221 33 -187
rect -33 -255 33 -221
rect -33 -289 -17 -255
rect 17 -289 33 -255
rect -33 -323 33 -289
rect -33 -357 -17 -323
rect 17 -357 33 -323
rect -33 -391 33 -357
rect -33 -425 -17 -391
rect 17 -425 33 -391
rect -33 -459 33 -425
rect -33 -493 -17 -459
rect 17 -493 33 -459
rect -33 -527 33 -493
rect -33 -561 -17 -527
rect 17 -561 33 -527
rect -33 -595 33 -561
rect -33 -629 -17 -595
rect 17 -629 33 -595
rect -33 -663 33 -629
rect -33 -697 -17 -663
rect 17 -697 33 -663
rect -33 -731 33 -697
rect -33 -765 -17 -731
rect 17 -765 33 -731
rect -33 -799 33 -765
rect -33 -833 -17 -799
rect 17 -833 33 -799
rect -33 -867 33 -833
rect -33 -901 -17 -867
rect 17 -901 33 -867
rect -33 -935 33 -901
rect -33 -969 -17 -935
rect 17 -969 33 -935
rect -33 -1000 33 -969
rect 63 969 125 1000
rect 63 935 79 969
rect 113 935 125 969
rect 63 901 125 935
rect 63 867 79 901
rect 113 867 125 901
rect 63 833 125 867
rect 63 799 79 833
rect 113 799 125 833
rect 63 765 125 799
rect 63 731 79 765
rect 113 731 125 765
rect 63 697 125 731
rect 63 663 79 697
rect 113 663 125 697
rect 63 629 125 663
rect 63 595 79 629
rect 113 595 125 629
rect 63 561 125 595
rect 63 527 79 561
rect 113 527 125 561
rect 63 493 125 527
rect 63 459 79 493
rect 113 459 125 493
rect 63 425 125 459
rect 63 391 79 425
rect 113 391 125 425
rect 63 357 125 391
rect 63 323 79 357
rect 113 323 125 357
rect 63 289 125 323
rect 63 255 79 289
rect 113 255 125 289
rect 63 221 125 255
rect 63 187 79 221
rect 113 187 125 221
rect 63 153 125 187
rect 63 119 79 153
rect 113 119 125 153
rect 63 85 125 119
rect 63 51 79 85
rect 113 51 125 85
rect 63 17 125 51
rect 63 -17 79 17
rect 113 -17 125 17
rect 63 -51 125 -17
rect 63 -85 79 -51
rect 113 -85 125 -51
rect 63 -119 125 -85
rect 63 -153 79 -119
rect 113 -153 125 -119
rect 63 -187 125 -153
rect 63 -221 79 -187
rect 113 -221 125 -187
rect 63 -255 125 -221
rect 63 -289 79 -255
rect 113 -289 125 -255
rect 63 -323 125 -289
rect 63 -357 79 -323
rect 113 -357 125 -323
rect 63 -391 125 -357
rect 63 -425 79 -391
rect 113 -425 125 -391
rect 63 -459 125 -425
rect 63 -493 79 -459
rect 113 -493 125 -459
rect 63 -527 125 -493
rect 63 -561 79 -527
rect 113 -561 125 -527
rect 63 -595 125 -561
rect 63 -629 79 -595
rect 113 -629 125 -595
rect 63 -663 125 -629
rect 63 -697 79 -663
rect 113 -697 125 -663
rect 63 -731 125 -697
rect 63 -765 79 -731
rect 113 -765 125 -731
rect 63 -799 125 -765
rect 63 -833 79 -799
rect 113 -833 125 -799
rect 63 -867 125 -833
rect 63 -901 79 -867
rect 113 -901 125 -867
rect 63 -935 125 -901
rect 63 -969 79 -935
rect 113 -969 125 -935
rect 63 -1000 125 -969
<< pdiffc >>
rect -113 935 -79 969
rect -113 867 -79 901
rect -113 799 -79 833
rect -113 731 -79 765
rect -113 663 -79 697
rect -113 595 -79 629
rect -113 527 -79 561
rect -113 459 -79 493
rect -113 391 -79 425
rect -113 323 -79 357
rect -113 255 -79 289
rect -113 187 -79 221
rect -113 119 -79 153
rect -113 51 -79 85
rect -113 -17 -79 17
rect -113 -85 -79 -51
rect -113 -153 -79 -119
rect -113 -221 -79 -187
rect -113 -289 -79 -255
rect -113 -357 -79 -323
rect -113 -425 -79 -391
rect -113 -493 -79 -459
rect -113 -561 -79 -527
rect -113 -629 -79 -595
rect -113 -697 -79 -663
rect -113 -765 -79 -731
rect -113 -833 -79 -799
rect -113 -901 -79 -867
rect -113 -969 -79 -935
rect -17 935 17 969
rect -17 867 17 901
rect -17 799 17 833
rect -17 731 17 765
rect -17 663 17 697
rect -17 595 17 629
rect -17 527 17 561
rect -17 459 17 493
rect -17 391 17 425
rect -17 323 17 357
rect -17 255 17 289
rect -17 187 17 221
rect -17 119 17 153
rect -17 51 17 85
rect -17 -17 17 17
rect -17 -85 17 -51
rect -17 -153 17 -119
rect -17 -221 17 -187
rect -17 -289 17 -255
rect -17 -357 17 -323
rect -17 -425 17 -391
rect -17 -493 17 -459
rect -17 -561 17 -527
rect -17 -629 17 -595
rect -17 -697 17 -663
rect -17 -765 17 -731
rect -17 -833 17 -799
rect -17 -901 17 -867
rect -17 -969 17 -935
rect 79 935 113 969
rect 79 867 113 901
rect 79 799 113 833
rect 79 731 113 765
rect 79 663 113 697
rect 79 595 113 629
rect 79 527 113 561
rect 79 459 113 493
rect 79 391 113 425
rect 79 323 113 357
rect 79 255 113 289
rect 79 187 113 221
rect 79 119 113 153
rect 79 51 113 85
rect 79 -17 113 17
rect 79 -85 113 -51
rect 79 -153 113 -119
rect 79 -221 113 -187
rect 79 -289 113 -255
rect 79 -357 113 -323
rect 79 -425 113 -391
rect 79 -493 113 -459
rect 79 -561 113 -527
rect 79 -629 113 -595
rect 79 -697 113 -663
rect 79 -765 113 -731
rect 79 -833 113 -799
rect 79 -901 113 -867
rect 79 -969 113 -935
<< poly >>
rect -63 1000 -33 1026
rect 33 1000 63 1026
rect -63 -1026 -33 -1000
rect 33 -1026 63 -1000
rect -63 -1056 63 -1026
<< locali >>
rect -113 969 -79 1004
rect -113 901 -79 919
rect -113 833 -79 847
rect -113 765 -79 775
rect -113 697 -79 703
rect -113 629 -79 631
rect -113 593 -79 595
rect -113 521 -79 527
rect -113 449 -79 459
rect -113 377 -79 391
rect -113 305 -79 323
rect -113 233 -79 255
rect -113 161 -79 187
rect -113 89 -79 119
rect -113 17 -79 51
rect -113 -51 -79 -17
rect -113 -119 -79 -89
rect -113 -187 -79 -161
rect -113 -255 -79 -233
rect -113 -323 -79 -305
rect -113 -391 -79 -377
rect -113 -459 -79 -449
rect -113 -527 -79 -521
rect -113 -595 -79 -593
rect -113 -631 -79 -629
rect -113 -703 -79 -697
rect -113 -775 -79 -765
rect -113 -847 -79 -833
rect -113 -919 -79 -901
rect -113 -1004 -79 -969
rect -17 969 17 1004
rect -17 901 17 919
rect -17 833 17 847
rect -17 765 17 775
rect -17 697 17 703
rect -17 629 17 631
rect -17 593 17 595
rect -17 521 17 527
rect -17 449 17 459
rect -17 377 17 391
rect -17 305 17 323
rect -17 233 17 255
rect -17 161 17 187
rect -17 89 17 119
rect -17 17 17 51
rect -17 -51 17 -17
rect -17 -119 17 -89
rect -17 -187 17 -161
rect -17 -255 17 -233
rect -17 -323 17 -305
rect -17 -391 17 -377
rect -17 -459 17 -449
rect -17 -527 17 -521
rect -17 -595 17 -593
rect -17 -631 17 -629
rect -17 -703 17 -697
rect -17 -775 17 -765
rect -17 -847 17 -833
rect -17 -919 17 -901
rect -17 -1004 17 -969
rect 79 969 113 1004
rect 79 901 113 919
rect 79 833 113 847
rect 79 765 113 775
rect 79 697 113 703
rect 79 629 113 631
rect 79 593 113 595
rect 79 521 113 527
rect 79 449 113 459
rect 79 377 113 391
rect 79 305 113 323
rect 79 233 113 255
rect 79 161 113 187
rect 79 89 113 119
rect 79 17 113 51
rect 79 -51 113 -17
rect 79 -119 113 -89
rect 79 -187 113 -161
rect 79 -255 113 -233
rect 79 -323 113 -305
rect 79 -391 113 -377
rect 79 -459 113 -449
rect 79 -527 113 -521
rect 79 -595 113 -593
rect 79 -631 113 -629
rect 79 -703 113 -697
rect 79 -775 113 -765
rect 79 -847 113 -833
rect 79 -919 113 -901
rect 79 -1004 113 -969
<< viali >>
rect -113 935 -79 953
rect -113 919 -79 935
rect -113 867 -79 881
rect -113 847 -79 867
rect -113 799 -79 809
rect -113 775 -79 799
rect -113 731 -79 737
rect -113 703 -79 731
rect -113 663 -79 665
rect -113 631 -79 663
rect -113 561 -79 593
rect -113 559 -79 561
rect -113 493 -79 521
rect -113 487 -79 493
rect -113 425 -79 449
rect -113 415 -79 425
rect -113 357 -79 377
rect -113 343 -79 357
rect -113 289 -79 305
rect -113 271 -79 289
rect -113 221 -79 233
rect -113 199 -79 221
rect -113 153 -79 161
rect -113 127 -79 153
rect -113 85 -79 89
rect -113 55 -79 85
rect -113 -17 -79 17
rect -113 -85 -79 -55
rect -113 -89 -79 -85
rect -113 -153 -79 -127
rect -113 -161 -79 -153
rect -113 -221 -79 -199
rect -113 -233 -79 -221
rect -113 -289 -79 -271
rect -113 -305 -79 -289
rect -113 -357 -79 -343
rect -113 -377 -79 -357
rect -113 -425 -79 -415
rect -113 -449 -79 -425
rect -113 -493 -79 -487
rect -113 -521 -79 -493
rect -113 -561 -79 -559
rect -113 -593 -79 -561
rect -113 -663 -79 -631
rect -113 -665 -79 -663
rect -113 -731 -79 -703
rect -113 -737 -79 -731
rect -113 -799 -79 -775
rect -113 -809 -79 -799
rect -113 -867 -79 -847
rect -113 -881 -79 -867
rect -113 -935 -79 -919
rect -113 -953 -79 -935
rect -17 935 17 953
rect -17 919 17 935
rect -17 867 17 881
rect -17 847 17 867
rect -17 799 17 809
rect -17 775 17 799
rect -17 731 17 737
rect -17 703 17 731
rect -17 663 17 665
rect -17 631 17 663
rect -17 561 17 593
rect -17 559 17 561
rect -17 493 17 521
rect -17 487 17 493
rect -17 425 17 449
rect -17 415 17 425
rect -17 357 17 377
rect -17 343 17 357
rect -17 289 17 305
rect -17 271 17 289
rect -17 221 17 233
rect -17 199 17 221
rect -17 153 17 161
rect -17 127 17 153
rect -17 85 17 89
rect -17 55 17 85
rect -17 -17 17 17
rect -17 -85 17 -55
rect -17 -89 17 -85
rect -17 -153 17 -127
rect -17 -161 17 -153
rect -17 -221 17 -199
rect -17 -233 17 -221
rect -17 -289 17 -271
rect -17 -305 17 -289
rect -17 -357 17 -343
rect -17 -377 17 -357
rect -17 -425 17 -415
rect -17 -449 17 -425
rect -17 -493 17 -487
rect -17 -521 17 -493
rect -17 -561 17 -559
rect -17 -593 17 -561
rect -17 -663 17 -631
rect -17 -665 17 -663
rect -17 -731 17 -703
rect -17 -737 17 -731
rect -17 -799 17 -775
rect -17 -809 17 -799
rect -17 -867 17 -847
rect -17 -881 17 -867
rect -17 -935 17 -919
rect -17 -953 17 -935
rect 79 935 113 953
rect 79 919 113 935
rect 79 867 113 881
rect 79 847 113 867
rect 79 799 113 809
rect 79 775 113 799
rect 79 731 113 737
rect 79 703 113 731
rect 79 663 113 665
rect 79 631 113 663
rect 79 561 113 593
rect 79 559 113 561
rect 79 493 113 521
rect 79 487 113 493
rect 79 425 113 449
rect 79 415 113 425
rect 79 357 113 377
rect 79 343 113 357
rect 79 289 113 305
rect 79 271 113 289
rect 79 221 113 233
rect 79 199 113 221
rect 79 153 113 161
rect 79 127 113 153
rect 79 85 113 89
rect 79 55 113 85
rect 79 -17 113 17
rect 79 -85 113 -55
rect 79 -89 113 -85
rect 79 -153 113 -127
rect 79 -161 113 -153
rect 79 -221 113 -199
rect 79 -233 113 -221
rect 79 -289 113 -271
rect 79 -305 113 -289
rect 79 -357 113 -343
rect 79 -377 113 -357
rect 79 -425 113 -415
rect 79 -449 113 -425
rect 79 -493 113 -487
rect 79 -521 113 -493
rect 79 -561 113 -559
rect 79 -593 113 -561
rect 79 -663 113 -631
rect 79 -665 113 -663
rect 79 -731 113 -703
rect 79 -737 113 -731
rect 79 -799 113 -775
rect 79 -809 113 -799
rect 79 -867 113 -847
rect 79 -881 113 -867
rect 79 -935 113 -919
rect 79 -953 113 -935
<< metal1 >>
rect -119 953 -73 1000
rect -119 919 -113 953
rect -79 919 -73 953
rect -119 881 -73 919
rect -119 847 -113 881
rect -79 847 -73 881
rect -119 809 -73 847
rect -119 775 -113 809
rect -79 775 -73 809
rect -119 737 -73 775
rect -119 703 -113 737
rect -79 703 -73 737
rect -119 665 -73 703
rect -119 631 -113 665
rect -79 631 -73 665
rect -119 593 -73 631
rect -119 559 -113 593
rect -79 559 -73 593
rect -119 521 -73 559
rect -119 487 -113 521
rect -79 487 -73 521
rect -119 449 -73 487
rect -119 415 -113 449
rect -79 415 -73 449
rect -119 377 -73 415
rect -119 343 -113 377
rect -79 343 -73 377
rect -119 305 -73 343
rect -119 271 -113 305
rect -79 271 -73 305
rect -119 233 -73 271
rect -119 199 -113 233
rect -79 199 -73 233
rect -119 161 -73 199
rect -119 127 -113 161
rect -79 127 -73 161
rect -119 89 -73 127
rect -119 55 -113 89
rect -79 55 -73 89
rect -119 17 -73 55
rect -119 -17 -113 17
rect -79 -17 -73 17
rect -119 -55 -73 -17
rect -119 -89 -113 -55
rect -79 -89 -73 -55
rect -119 -127 -73 -89
rect -119 -161 -113 -127
rect -79 -161 -73 -127
rect -119 -199 -73 -161
rect -119 -233 -113 -199
rect -79 -233 -73 -199
rect -119 -271 -73 -233
rect -119 -305 -113 -271
rect -79 -305 -73 -271
rect -119 -343 -73 -305
rect -119 -377 -113 -343
rect -79 -377 -73 -343
rect -119 -415 -73 -377
rect -119 -449 -113 -415
rect -79 -449 -73 -415
rect -119 -487 -73 -449
rect -119 -521 -113 -487
rect -79 -521 -73 -487
rect -119 -559 -73 -521
rect -119 -593 -113 -559
rect -79 -593 -73 -559
rect -119 -631 -73 -593
rect -119 -665 -113 -631
rect -79 -665 -73 -631
rect -119 -703 -73 -665
rect -119 -737 -113 -703
rect -79 -737 -73 -703
rect -119 -775 -73 -737
rect -119 -809 -113 -775
rect -79 -809 -73 -775
rect -119 -847 -73 -809
rect -119 -881 -113 -847
rect -79 -881 -73 -847
rect -119 -919 -73 -881
rect -119 -953 -113 -919
rect -79 -953 -73 -919
rect -119 -1000 -73 -953
rect -23 953 23 1000
rect -23 919 -17 953
rect 17 919 23 953
rect -23 881 23 919
rect -23 847 -17 881
rect 17 847 23 881
rect -23 809 23 847
rect -23 775 -17 809
rect 17 775 23 809
rect -23 737 23 775
rect -23 703 -17 737
rect 17 703 23 737
rect -23 665 23 703
rect -23 631 -17 665
rect 17 631 23 665
rect -23 593 23 631
rect -23 559 -17 593
rect 17 559 23 593
rect -23 521 23 559
rect -23 487 -17 521
rect 17 487 23 521
rect -23 449 23 487
rect -23 415 -17 449
rect 17 415 23 449
rect -23 377 23 415
rect -23 343 -17 377
rect 17 343 23 377
rect -23 305 23 343
rect -23 271 -17 305
rect 17 271 23 305
rect -23 233 23 271
rect -23 199 -17 233
rect 17 199 23 233
rect -23 161 23 199
rect -23 127 -17 161
rect 17 127 23 161
rect -23 89 23 127
rect -23 55 -17 89
rect 17 55 23 89
rect -23 17 23 55
rect -23 -17 -17 17
rect 17 -17 23 17
rect -23 -55 23 -17
rect -23 -89 -17 -55
rect 17 -89 23 -55
rect -23 -127 23 -89
rect -23 -161 -17 -127
rect 17 -161 23 -127
rect -23 -199 23 -161
rect -23 -233 -17 -199
rect 17 -233 23 -199
rect -23 -271 23 -233
rect -23 -305 -17 -271
rect 17 -305 23 -271
rect -23 -343 23 -305
rect -23 -377 -17 -343
rect 17 -377 23 -343
rect -23 -415 23 -377
rect -23 -449 -17 -415
rect 17 -449 23 -415
rect -23 -487 23 -449
rect -23 -521 -17 -487
rect 17 -521 23 -487
rect -23 -559 23 -521
rect -23 -593 -17 -559
rect 17 -593 23 -559
rect -23 -631 23 -593
rect -23 -665 -17 -631
rect 17 -665 23 -631
rect -23 -703 23 -665
rect -23 -737 -17 -703
rect 17 -737 23 -703
rect -23 -775 23 -737
rect -23 -809 -17 -775
rect 17 -809 23 -775
rect -23 -847 23 -809
rect -23 -881 -17 -847
rect 17 -881 23 -847
rect -23 -919 23 -881
rect -23 -953 -17 -919
rect 17 -953 23 -919
rect -23 -1000 23 -953
rect 73 953 119 1000
rect 73 919 79 953
rect 113 919 119 953
rect 73 881 119 919
rect 73 847 79 881
rect 113 847 119 881
rect 73 809 119 847
rect 73 775 79 809
rect 113 775 119 809
rect 73 737 119 775
rect 73 703 79 737
rect 113 703 119 737
rect 73 665 119 703
rect 73 631 79 665
rect 113 631 119 665
rect 73 593 119 631
rect 73 559 79 593
rect 113 559 119 593
rect 73 521 119 559
rect 73 487 79 521
rect 113 487 119 521
rect 73 449 119 487
rect 73 415 79 449
rect 113 415 119 449
rect 73 377 119 415
rect 73 343 79 377
rect 113 343 119 377
rect 73 305 119 343
rect 73 271 79 305
rect 113 271 119 305
rect 73 233 119 271
rect 73 199 79 233
rect 113 199 119 233
rect 73 161 119 199
rect 73 127 79 161
rect 113 127 119 161
rect 73 89 119 127
rect 73 55 79 89
rect 113 55 119 89
rect 73 17 119 55
rect 73 -17 79 17
rect 113 -17 119 17
rect 73 -55 119 -17
rect 73 -89 79 -55
rect 113 -89 119 -55
rect 73 -127 119 -89
rect 73 -161 79 -127
rect 113 -161 119 -127
rect 73 -199 119 -161
rect 73 -233 79 -199
rect 113 -233 119 -199
rect 73 -271 119 -233
rect 73 -305 79 -271
rect 113 -305 119 -271
rect 73 -343 119 -305
rect 73 -377 79 -343
rect 113 -377 119 -343
rect 73 -415 119 -377
rect 73 -449 79 -415
rect 113 -449 119 -415
rect 73 -487 119 -449
rect 73 -521 79 -487
rect 113 -521 119 -487
rect 73 -559 119 -521
rect 73 -593 79 -559
rect 113 -593 119 -559
rect 73 -631 119 -593
rect 73 -665 79 -631
rect 113 -665 119 -631
rect 73 -703 119 -665
rect 73 -737 79 -703
rect 113 -737 119 -703
rect 73 -775 119 -737
rect 73 -809 79 -775
rect 113 -809 119 -775
rect 73 -847 119 -809
rect 73 -881 79 -847
rect 113 -881 119 -847
rect 73 -919 119 -881
rect 73 -953 79 -919
rect 113 -953 119 -919
rect 73 -1000 119 -953
<< end >>
