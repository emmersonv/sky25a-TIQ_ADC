** sch_path: /foss/designs/analog-circuit-design/sky25a-TIQ_ADC/xschem/gain_stage.sch
.subckt gain_stage in out VGND VDPWR
*.PININFO in:I out:O VGND:B VDPWR:B
x8 VDPWR net1 in VGND inverter_p1_n0o42
x9 VDPWR net2 net1 VGND inverter_p1_n0o42
x10 VDPWR out net2 VGND inverter_p1_n0o42
.ends

* expanding   symbol:  /foss/designs/analog-circuit-design/sky25a-TIQ_ADC/xschem/INVERTER_SIZES/inverter_p1_n0o42.sym # of pins=4
** sym_path: /foss/designs/analog-circuit-design/sky25a-TIQ_ADC/xschem/INVERTER_SIZES/inverter_p1_n0o42.sym
** sch_path: /foss/designs/analog-circuit-design/sky25a-TIQ_ADC/xschem/INVERTER_SIZES/inverter_p1_n0o42.sch
.subckt inverter_p1_n0o42 VDPWR Vout Vin VGND
*.PININFO Vout:O Vin:I VDPWR:B VGND:B
XM1 Vout Vin VGND VGND sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM2 Vout Vin VDPWR VDPWR sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 m=1
.ends

