magic
tech sky130A
magscale 1 2
timestamp 1756008383
<< nwell >>
rect -209 -1062 209 1062
<< pmos >>
rect -111 -1000 -81 1000
rect -15 -1000 15 1000
rect 81 -1000 111 1000
<< pdiff >>
rect -173 969 -111 1000
rect -173 935 -161 969
rect -127 935 -111 969
rect -173 901 -111 935
rect -173 867 -161 901
rect -127 867 -111 901
rect -173 833 -111 867
rect -173 799 -161 833
rect -127 799 -111 833
rect -173 765 -111 799
rect -173 731 -161 765
rect -127 731 -111 765
rect -173 697 -111 731
rect -173 663 -161 697
rect -127 663 -111 697
rect -173 629 -111 663
rect -173 595 -161 629
rect -127 595 -111 629
rect -173 561 -111 595
rect -173 527 -161 561
rect -127 527 -111 561
rect -173 493 -111 527
rect -173 459 -161 493
rect -127 459 -111 493
rect -173 425 -111 459
rect -173 391 -161 425
rect -127 391 -111 425
rect -173 357 -111 391
rect -173 323 -161 357
rect -127 323 -111 357
rect -173 289 -111 323
rect -173 255 -161 289
rect -127 255 -111 289
rect -173 221 -111 255
rect -173 187 -161 221
rect -127 187 -111 221
rect -173 153 -111 187
rect -173 119 -161 153
rect -127 119 -111 153
rect -173 85 -111 119
rect -173 51 -161 85
rect -127 51 -111 85
rect -173 17 -111 51
rect -173 -17 -161 17
rect -127 -17 -111 17
rect -173 -51 -111 -17
rect -173 -85 -161 -51
rect -127 -85 -111 -51
rect -173 -119 -111 -85
rect -173 -153 -161 -119
rect -127 -153 -111 -119
rect -173 -187 -111 -153
rect -173 -221 -161 -187
rect -127 -221 -111 -187
rect -173 -255 -111 -221
rect -173 -289 -161 -255
rect -127 -289 -111 -255
rect -173 -323 -111 -289
rect -173 -357 -161 -323
rect -127 -357 -111 -323
rect -173 -391 -111 -357
rect -173 -425 -161 -391
rect -127 -425 -111 -391
rect -173 -459 -111 -425
rect -173 -493 -161 -459
rect -127 -493 -111 -459
rect -173 -527 -111 -493
rect -173 -561 -161 -527
rect -127 -561 -111 -527
rect -173 -595 -111 -561
rect -173 -629 -161 -595
rect -127 -629 -111 -595
rect -173 -663 -111 -629
rect -173 -697 -161 -663
rect -127 -697 -111 -663
rect -173 -731 -111 -697
rect -173 -765 -161 -731
rect -127 -765 -111 -731
rect -173 -799 -111 -765
rect -173 -833 -161 -799
rect -127 -833 -111 -799
rect -173 -867 -111 -833
rect -173 -901 -161 -867
rect -127 -901 -111 -867
rect -173 -935 -111 -901
rect -173 -969 -161 -935
rect -127 -969 -111 -935
rect -173 -1000 -111 -969
rect -81 969 -15 1000
rect -81 935 -65 969
rect -31 935 -15 969
rect -81 901 -15 935
rect -81 867 -65 901
rect -31 867 -15 901
rect -81 833 -15 867
rect -81 799 -65 833
rect -31 799 -15 833
rect -81 765 -15 799
rect -81 731 -65 765
rect -31 731 -15 765
rect -81 697 -15 731
rect -81 663 -65 697
rect -31 663 -15 697
rect -81 629 -15 663
rect -81 595 -65 629
rect -31 595 -15 629
rect -81 561 -15 595
rect -81 527 -65 561
rect -31 527 -15 561
rect -81 493 -15 527
rect -81 459 -65 493
rect -31 459 -15 493
rect -81 425 -15 459
rect -81 391 -65 425
rect -31 391 -15 425
rect -81 357 -15 391
rect -81 323 -65 357
rect -31 323 -15 357
rect -81 289 -15 323
rect -81 255 -65 289
rect -31 255 -15 289
rect -81 221 -15 255
rect -81 187 -65 221
rect -31 187 -15 221
rect -81 153 -15 187
rect -81 119 -65 153
rect -31 119 -15 153
rect -81 85 -15 119
rect -81 51 -65 85
rect -31 51 -15 85
rect -81 17 -15 51
rect -81 -17 -65 17
rect -31 -17 -15 17
rect -81 -51 -15 -17
rect -81 -85 -65 -51
rect -31 -85 -15 -51
rect -81 -119 -15 -85
rect -81 -153 -65 -119
rect -31 -153 -15 -119
rect -81 -187 -15 -153
rect -81 -221 -65 -187
rect -31 -221 -15 -187
rect -81 -255 -15 -221
rect -81 -289 -65 -255
rect -31 -289 -15 -255
rect -81 -323 -15 -289
rect -81 -357 -65 -323
rect -31 -357 -15 -323
rect -81 -391 -15 -357
rect -81 -425 -65 -391
rect -31 -425 -15 -391
rect -81 -459 -15 -425
rect -81 -493 -65 -459
rect -31 -493 -15 -459
rect -81 -527 -15 -493
rect -81 -561 -65 -527
rect -31 -561 -15 -527
rect -81 -595 -15 -561
rect -81 -629 -65 -595
rect -31 -629 -15 -595
rect -81 -663 -15 -629
rect -81 -697 -65 -663
rect -31 -697 -15 -663
rect -81 -731 -15 -697
rect -81 -765 -65 -731
rect -31 -765 -15 -731
rect -81 -799 -15 -765
rect -81 -833 -65 -799
rect -31 -833 -15 -799
rect -81 -867 -15 -833
rect -81 -901 -65 -867
rect -31 -901 -15 -867
rect -81 -935 -15 -901
rect -81 -969 -65 -935
rect -31 -969 -15 -935
rect -81 -1000 -15 -969
rect 15 969 81 1000
rect 15 935 31 969
rect 65 935 81 969
rect 15 901 81 935
rect 15 867 31 901
rect 65 867 81 901
rect 15 833 81 867
rect 15 799 31 833
rect 65 799 81 833
rect 15 765 81 799
rect 15 731 31 765
rect 65 731 81 765
rect 15 697 81 731
rect 15 663 31 697
rect 65 663 81 697
rect 15 629 81 663
rect 15 595 31 629
rect 65 595 81 629
rect 15 561 81 595
rect 15 527 31 561
rect 65 527 81 561
rect 15 493 81 527
rect 15 459 31 493
rect 65 459 81 493
rect 15 425 81 459
rect 15 391 31 425
rect 65 391 81 425
rect 15 357 81 391
rect 15 323 31 357
rect 65 323 81 357
rect 15 289 81 323
rect 15 255 31 289
rect 65 255 81 289
rect 15 221 81 255
rect 15 187 31 221
rect 65 187 81 221
rect 15 153 81 187
rect 15 119 31 153
rect 65 119 81 153
rect 15 85 81 119
rect 15 51 31 85
rect 65 51 81 85
rect 15 17 81 51
rect 15 -17 31 17
rect 65 -17 81 17
rect 15 -51 81 -17
rect 15 -85 31 -51
rect 65 -85 81 -51
rect 15 -119 81 -85
rect 15 -153 31 -119
rect 65 -153 81 -119
rect 15 -187 81 -153
rect 15 -221 31 -187
rect 65 -221 81 -187
rect 15 -255 81 -221
rect 15 -289 31 -255
rect 65 -289 81 -255
rect 15 -323 81 -289
rect 15 -357 31 -323
rect 65 -357 81 -323
rect 15 -391 81 -357
rect 15 -425 31 -391
rect 65 -425 81 -391
rect 15 -459 81 -425
rect 15 -493 31 -459
rect 65 -493 81 -459
rect 15 -527 81 -493
rect 15 -561 31 -527
rect 65 -561 81 -527
rect 15 -595 81 -561
rect 15 -629 31 -595
rect 65 -629 81 -595
rect 15 -663 81 -629
rect 15 -697 31 -663
rect 65 -697 81 -663
rect 15 -731 81 -697
rect 15 -765 31 -731
rect 65 -765 81 -731
rect 15 -799 81 -765
rect 15 -833 31 -799
rect 65 -833 81 -799
rect 15 -867 81 -833
rect 15 -901 31 -867
rect 65 -901 81 -867
rect 15 -935 81 -901
rect 15 -969 31 -935
rect 65 -969 81 -935
rect 15 -1000 81 -969
rect 111 969 173 1000
rect 111 935 127 969
rect 161 935 173 969
rect 111 901 173 935
rect 111 867 127 901
rect 161 867 173 901
rect 111 833 173 867
rect 111 799 127 833
rect 161 799 173 833
rect 111 765 173 799
rect 111 731 127 765
rect 161 731 173 765
rect 111 697 173 731
rect 111 663 127 697
rect 161 663 173 697
rect 111 629 173 663
rect 111 595 127 629
rect 161 595 173 629
rect 111 561 173 595
rect 111 527 127 561
rect 161 527 173 561
rect 111 493 173 527
rect 111 459 127 493
rect 161 459 173 493
rect 111 425 173 459
rect 111 391 127 425
rect 161 391 173 425
rect 111 357 173 391
rect 111 323 127 357
rect 161 323 173 357
rect 111 289 173 323
rect 111 255 127 289
rect 161 255 173 289
rect 111 221 173 255
rect 111 187 127 221
rect 161 187 173 221
rect 111 153 173 187
rect 111 119 127 153
rect 161 119 173 153
rect 111 85 173 119
rect 111 51 127 85
rect 161 51 173 85
rect 111 17 173 51
rect 111 -17 127 17
rect 161 -17 173 17
rect 111 -51 173 -17
rect 111 -85 127 -51
rect 161 -85 173 -51
rect 111 -119 173 -85
rect 111 -153 127 -119
rect 161 -153 173 -119
rect 111 -187 173 -153
rect 111 -221 127 -187
rect 161 -221 173 -187
rect 111 -255 173 -221
rect 111 -289 127 -255
rect 161 -289 173 -255
rect 111 -323 173 -289
rect 111 -357 127 -323
rect 161 -357 173 -323
rect 111 -391 173 -357
rect 111 -425 127 -391
rect 161 -425 173 -391
rect 111 -459 173 -425
rect 111 -493 127 -459
rect 161 -493 173 -459
rect 111 -527 173 -493
rect 111 -561 127 -527
rect 161 -561 173 -527
rect 111 -595 173 -561
rect 111 -629 127 -595
rect 161 -629 173 -595
rect 111 -663 173 -629
rect 111 -697 127 -663
rect 161 -697 173 -663
rect 111 -731 173 -697
rect 111 -765 127 -731
rect 161 -765 173 -731
rect 111 -799 173 -765
rect 111 -833 127 -799
rect 161 -833 173 -799
rect 111 -867 173 -833
rect 111 -901 127 -867
rect 161 -901 173 -867
rect 111 -935 173 -901
rect 111 -969 127 -935
rect 161 -969 173 -935
rect 111 -1000 173 -969
<< pdiffc >>
rect -161 935 -127 969
rect -161 867 -127 901
rect -161 799 -127 833
rect -161 731 -127 765
rect -161 663 -127 697
rect -161 595 -127 629
rect -161 527 -127 561
rect -161 459 -127 493
rect -161 391 -127 425
rect -161 323 -127 357
rect -161 255 -127 289
rect -161 187 -127 221
rect -161 119 -127 153
rect -161 51 -127 85
rect -161 -17 -127 17
rect -161 -85 -127 -51
rect -161 -153 -127 -119
rect -161 -221 -127 -187
rect -161 -289 -127 -255
rect -161 -357 -127 -323
rect -161 -425 -127 -391
rect -161 -493 -127 -459
rect -161 -561 -127 -527
rect -161 -629 -127 -595
rect -161 -697 -127 -663
rect -161 -765 -127 -731
rect -161 -833 -127 -799
rect -161 -901 -127 -867
rect -161 -969 -127 -935
rect -65 935 -31 969
rect -65 867 -31 901
rect -65 799 -31 833
rect -65 731 -31 765
rect -65 663 -31 697
rect -65 595 -31 629
rect -65 527 -31 561
rect -65 459 -31 493
rect -65 391 -31 425
rect -65 323 -31 357
rect -65 255 -31 289
rect -65 187 -31 221
rect -65 119 -31 153
rect -65 51 -31 85
rect -65 -17 -31 17
rect -65 -85 -31 -51
rect -65 -153 -31 -119
rect -65 -221 -31 -187
rect -65 -289 -31 -255
rect -65 -357 -31 -323
rect -65 -425 -31 -391
rect -65 -493 -31 -459
rect -65 -561 -31 -527
rect -65 -629 -31 -595
rect -65 -697 -31 -663
rect -65 -765 -31 -731
rect -65 -833 -31 -799
rect -65 -901 -31 -867
rect -65 -969 -31 -935
rect 31 935 65 969
rect 31 867 65 901
rect 31 799 65 833
rect 31 731 65 765
rect 31 663 65 697
rect 31 595 65 629
rect 31 527 65 561
rect 31 459 65 493
rect 31 391 65 425
rect 31 323 65 357
rect 31 255 65 289
rect 31 187 65 221
rect 31 119 65 153
rect 31 51 65 85
rect 31 -17 65 17
rect 31 -85 65 -51
rect 31 -153 65 -119
rect 31 -221 65 -187
rect 31 -289 65 -255
rect 31 -357 65 -323
rect 31 -425 65 -391
rect 31 -493 65 -459
rect 31 -561 65 -527
rect 31 -629 65 -595
rect 31 -697 65 -663
rect 31 -765 65 -731
rect 31 -833 65 -799
rect 31 -901 65 -867
rect 31 -969 65 -935
rect 127 935 161 969
rect 127 867 161 901
rect 127 799 161 833
rect 127 731 161 765
rect 127 663 161 697
rect 127 595 161 629
rect 127 527 161 561
rect 127 459 161 493
rect 127 391 161 425
rect 127 323 161 357
rect 127 255 161 289
rect 127 187 161 221
rect 127 119 161 153
rect 127 51 161 85
rect 127 -17 161 17
rect 127 -85 161 -51
rect 127 -153 161 -119
rect 127 -221 161 -187
rect 127 -289 161 -255
rect 127 -357 161 -323
rect 127 -425 161 -391
rect 127 -493 161 -459
rect 127 -561 161 -527
rect 127 -629 161 -595
rect 127 -697 161 -663
rect 127 -765 161 -731
rect 127 -833 161 -799
rect 127 -901 161 -867
rect 127 -969 161 -935
<< poly >>
rect -111 1000 -81 1026
rect -15 1000 15 1026
rect 81 1000 111 1026
rect -111 -1026 -81 -1000
rect -15 -1026 15 -1000
rect 81 -1026 111 -1000
rect -111 -1056 111 -1026
<< locali >>
rect -161 969 -127 1004
rect -161 901 -127 919
rect -161 833 -127 847
rect -161 765 -127 775
rect -161 697 -127 703
rect -161 629 -127 631
rect -161 593 -127 595
rect -161 521 -127 527
rect -161 449 -127 459
rect -161 377 -127 391
rect -161 305 -127 323
rect -161 233 -127 255
rect -161 161 -127 187
rect -161 89 -127 119
rect -161 17 -127 51
rect -161 -51 -127 -17
rect -161 -119 -127 -89
rect -161 -187 -127 -161
rect -161 -255 -127 -233
rect -161 -323 -127 -305
rect -161 -391 -127 -377
rect -161 -459 -127 -449
rect -161 -527 -127 -521
rect -161 -595 -127 -593
rect -161 -631 -127 -629
rect -161 -703 -127 -697
rect -161 -775 -127 -765
rect -161 -847 -127 -833
rect -161 -919 -127 -901
rect -161 -1004 -127 -969
rect -65 969 -31 1004
rect -65 901 -31 919
rect -65 833 -31 847
rect -65 765 -31 775
rect -65 697 -31 703
rect -65 629 -31 631
rect -65 593 -31 595
rect -65 521 -31 527
rect -65 449 -31 459
rect -65 377 -31 391
rect -65 305 -31 323
rect -65 233 -31 255
rect -65 161 -31 187
rect -65 89 -31 119
rect -65 17 -31 51
rect -65 -51 -31 -17
rect -65 -119 -31 -89
rect -65 -187 -31 -161
rect -65 -255 -31 -233
rect -65 -323 -31 -305
rect -65 -391 -31 -377
rect -65 -459 -31 -449
rect -65 -527 -31 -521
rect -65 -595 -31 -593
rect -65 -631 -31 -629
rect -65 -703 -31 -697
rect -65 -775 -31 -765
rect -65 -847 -31 -833
rect -65 -919 -31 -901
rect -65 -1004 -31 -969
rect 31 969 65 1004
rect 31 901 65 919
rect 31 833 65 847
rect 31 765 65 775
rect 31 697 65 703
rect 31 629 65 631
rect 31 593 65 595
rect 31 521 65 527
rect 31 449 65 459
rect 31 377 65 391
rect 31 305 65 323
rect 31 233 65 255
rect 31 161 65 187
rect 31 89 65 119
rect 31 17 65 51
rect 31 -51 65 -17
rect 31 -119 65 -89
rect 31 -187 65 -161
rect 31 -255 65 -233
rect 31 -323 65 -305
rect 31 -391 65 -377
rect 31 -459 65 -449
rect 31 -527 65 -521
rect 31 -595 65 -593
rect 31 -631 65 -629
rect 31 -703 65 -697
rect 31 -775 65 -765
rect 31 -847 65 -833
rect 31 -919 65 -901
rect 31 -1004 65 -969
rect 127 969 161 1004
rect 127 901 161 919
rect 127 833 161 847
rect 127 765 161 775
rect 127 697 161 703
rect 127 629 161 631
rect 127 593 161 595
rect 127 521 161 527
rect 127 449 161 459
rect 127 377 161 391
rect 127 305 161 323
rect 127 233 161 255
rect 127 161 161 187
rect 127 89 161 119
rect 127 17 161 51
rect 127 -51 161 -17
rect 127 -119 161 -89
rect 127 -187 161 -161
rect 127 -255 161 -233
rect 127 -323 161 -305
rect 127 -391 161 -377
rect 127 -459 161 -449
rect 127 -527 161 -521
rect 127 -595 161 -593
rect 127 -631 161 -629
rect 127 -703 161 -697
rect 127 -775 161 -765
rect 127 -847 161 -833
rect 127 -919 161 -901
rect 127 -1004 161 -969
<< viali >>
rect -161 935 -127 953
rect -161 919 -127 935
rect -161 867 -127 881
rect -161 847 -127 867
rect -161 799 -127 809
rect -161 775 -127 799
rect -161 731 -127 737
rect -161 703 -127 731
rect -161 663 -127 665
rect -161 631 -127 663
rect -161 561 -127 593
rect -161 559 -127 561
rect -161 493 -127 521
rect -161 487 -127 493
rect -161 425 -127 449
rect -161 415 -127 425
rect -161 357 -127 377
rect -161 343 -127 357
rect -161 289 -127 305
rect -161 271 -127 289
rect -161 221 -127 233
rect -161 199 -127 221
rect -161 153 -127 161
rect -161 127 -127 153
rect -161 85 -127 89
rect -161 55 -127 85
rect -161 -17 -127 17
rect -161 -85 -127 -55
rect -161 -89 -127 -85
rect -161 -153 -127 -127
rect -161 -161 -127 -153
rect -161 -221 -127 -199
rect -161 -233 -127 -221
rect -161 -289 -127 -271
rect -161 -305 -127 -289
rect -161 -357 -127 -343
rect -161 -377 -127 -357
rect -161 -425 -127 -415
rect -161 -449 -127 -425
rect -161 -493 -127 -487
rect -161 -521 -127 -493
rect -161 -561 -127 -559
rect -161 -593 -127 -561
rect -161 -663 -127 -631
rect -161 -665 -127 -663
rect -161 -731 -127 -703
rect -161 -737 -127 -731
rect -161 -799 -127 -775
rect -161 -809 -127 -799
rect -161 -867 -127 -847
rect -161 -881 -127 -867
rect -161 -935 -127 -919
rect -161 -953 -127 -935
rect -65 935 -31 953
rect -65 919 -31 935
rect -65 867 -31 881
rect -65 847 -31 867
rect -65 799 -31 809
rect -65 775 -31 799
rect -65 731 -31 737
rect -65 703 -31 731
rect -65 663 -31 665
rect -65 631 -31 663
rect -65 561 -31 593
rect -65 559 -31 561
rect -65 493 -31 521
rect -65 487 -31 493
rect -65 425 -31 449
rect -65 415 -31 425
rect -65 357 -31 377
rect -65 343 -31 357
rect -65 289 -31 305
rect -65 271 -31 289
rect -65 221 -31 233
rect -65 199 -31 221
rect -65 153 -31 161
rect -65 127 -31 153
rect -65 85 -31 89
rect -65 55 -31 85
rect -65 -17 -31 17
rect -65 -85 -31 -55
rect -65 -89 -31 -85
rect -65 -153 -31 -127
rect -65 -161 -31 -153
rect -65 -221 -31 -199
rect -65 -233 -31 -221
rect -65 -289 -31 -271
rect -65 -305 -31 -289
rect -65 -357 -31 -343
rect -65 -377 -31 -357
rect -65 -425 -31 -415
rect -65 -449 -31 -425
rect -65 -493 -31 -487
rect -65 -521 -31 -493
rect -65 -561 -31 -559
rect -65 -593 -31 -561
rect -65 -663 -31 -631
rect -65 -665 -31 -663
rect -65 -731 -31 -703
rect -65 -737 -31 -731
rect -65 -799 -31 -775
rect -65 -809 -31 -799
rect -65 -867 -31 -847
rect -65 -881 -31 -867
rect -65 -935 -31 -919
rect -65 -953 -31 -935
rect 31 935 65 953
rect 31 919 65 935
rect 31 867 65 881
rect 31 847 65 867
rect 31 799 65 809
rect 31 775 65 799
rect 31 731 65 737
rect 31 703 65 731
rect 31 663 65 665
rect 31 631 65 663
rect 31 561 65 593
rect 31 559 65 561
rect 31 493 65 521
rect 31 487 65 493
rect 31 425 65 449
rect 31 415 65 425
rect 31 357 65 377
rect 31 343 65 357
rect 31 289 65 305
rect 31 271 65 289
rect 31 221 65 233
rect 31 199 65 221
rect 31 153 65 161
rect 31 127 65 153
rect 31 85 65 89
rect 31 55 65 85
rect 31 -17 65 17
rect 31 -85 65 -55
rect 31 -89 65 -85
rect 31 -153 65 -127
rect 31 -161 65 -153
rect 31 -221 65 -199
rect 31 -233 65 -221
rect 31 -289 65 -271
rect 31 -305 65 -289
rect 31 -357 65 -343
rect 31 -377 65 -357
rect 31 -425 65 -415
rect 31 -449 65 -425
rect 31 -493 65 -487
rect 31 -521 65 -493
rect 31 -561 65 -559
rect 31 -593 65 -561
rect 31 -663 65 -631
rect 31 -665 65 -663
rect 31 -731 65 -703
rect 31 -737 65 -731
rect 31 -799 65 -775
rect 31 -809 65 -799
rect 31 -867 65 -847
rect 31 -881 65 -867
rect 31 -935 65 -919
rect 31 -953 65 -935
rect 127 935 161 953
rect 127 919 161 935
rect 127 867 161 881
rect 127 847 161 867
rect 127 799 161 809
rect 127 775 161 799
rect 127 731 161 737
rect 127 703 161 731
rect 127 663 161 665
rect 127 631 161 663
rect 127 561 161 593
rect 127 559 161 561
rect 127 493 161 521
rect 127 487 161 493
rect 127 425 161 449
rect 127 415 161 425
rect 127 357 161 377
rect 127 343 161 357
rect 127 289 161 305
rect 127 271 161 289
rect 127 221 161 233
rect 127 199 161 221
rect 127 153 161 161
rect 127 127 161 153
rect 127 85 161 89
rect 127 55 161 85
rect 127 -17 161 17
rect 127 -85 161 -55
rect 127 -89 161 -85
rect 127 -153 161 -127
rect 127 -161 161 -153
rect 127 -221 161 -199
rect 127 -233 161 -221
rect 127 -289 161 -271
rect 127 -305 161 -289
rect 127 -357 161 -343
rect 127 -377 161 -357
rect 127 -425 161 -415
rect 127 -449 161 -425
rect 127 -493 161 -487
rect 127 -521 161 -493
rect 127 -561 161 -559
rect 127 -593 161 -561
rect 127 -663 161 -631
rect 127 -665 161 -663
rect 127 -731 161 -703
rect 127 -737 161 -731
rect 127 -799 161 -775
rect 127 -809 161 -799
rect 127 -867 161 -847
rect 127 -881 161 -867
rect 127 -935 161 -919
rect 127 -953 161 -935
<< metal1 >>
rect -167 953 -121 1000
rect -167 919 -161 953
rect -127 919 -121 953
rect -167 881 -121 919
rect -167 847 -161 881
rect -127 847 -121 881
rect -167 809 -121 847
rect -167 775 -161 809
rect -127 775 -121 809
rect -167 737 -121 775
rect -167 703 -161 737
rect -127 703 -121 737
rect -167 665 -121 703
rect -167 631 -161 665
rect -127 631 -121 665
rect -167 593 -121 631
rect -167 559 -161 593
rect -127 559 -121 593
rect -167 521 -121 559
rect -167 487 -161 521
rect -127 487 -121 521
rect -167 449 -121 487
rect -167 415 -161 449
rect -127 415 -121 449
rect -167 377 -121 415
rect -167 343 -161 377
rect -127 343 -121 377
rect -167 305 -121 343
rect -167 271 -161 305
rect -127 271 -121 305
rect -167 233 -121 271
rect -167 199 -161 233
rect -127 199 -121 233
rect -167 161 -121 199
rect -167 127 -161 161
rect -127 127 -121 161
rect -167 89 -121 127
rect -167 55 -161 89
rect -127 55 -121 89
rect -167 17 -121 55
rect -167 -17 -161 17
rect -127 -17 -121 17
rect -167 -55 -121 -17
rect -167 -89 -161 -55
rect -127 -89 -121 -55
rect -167 -127 -121 -89
rect -167 -161 -161 -127
rect -127 -161 -121 -127
rect -167 -199 -121 -161
rect -167 -233 -161 -199
rect -127 -233 -121 -199
rect -167 -271 -121 -233
rect -167 -305 -161 -271
rect -127 -305 -121 -271
rect -167 -343 -121 -305
rect -167 -377 -161 -343
rect -127 -377 -121 -343
rect -167 -415 -121 -377
rect -167 -449 -161 -415
rect -127 -449 -121 -415
rect -167 -487 -121 -449
rect -167 -521 -161 -487
rect -127 -521 -121 -487
rect -167 -559 -121 -521
rect -167 -593 -161 -559
rect -127 -593 -121 -559
rect -167 -631 -121 -593
rect -167 -665 -161 -631
rect -127 -665 -121 -631
rect -167 -703 -121 -665
rect -167 -737 -161 -703
rect -127 -737 -121 -703
rect -167 -775 -121 -737
rect -167 -809 -161 -775
rect -127 -809 -121 -775
rect -167 -847 -121 -809
rect -167 -881 -161 -847
rect -127 -881 -121 -847
rect -167 -919 -121 -881
rect -167 -953 -161 -919
rect -127 -953 -121 -919
rect -167 -1000 -121 -953
rect -71 953 -25 1000
rect -71 919 -65 953
rect -31 919 -25 953
rect -71 881 -25 919
rect -71 847 -65 881
rect -31 847 -25 881
rect -71 809 -25 847
rect -71 775 -65 809
rect -31 775 -25 809
rect -71 737 -25 775
rect -71 703 -65 737
rect -31 703 -25 737
rect -71 665 -25 703
rect -71 631 -65 665
rect -31 631 -25 665
rect -71 593 -25 631
rect -71 559 -65 593
rect -31 559 -25 593
rect -71 521 -25 559
rect -71 487 -65 521
rect -31 487 -25 521
rect -71 449 -25 487
rect -71 415 -65 449
rect -31 415 -25 449
rect -71 377 -25 415
rect -71 343 -65 377
rect -31 343 -25 377
rect -71 305 -25 343
rect -71 271 -65 305
rect -31 271 -25 305
rect -71 233 -25 271
rect -71 199 -65 233
rect -31 199 -25 233
rect -71 161 -25 199
rect -71 127 -65 161
rect -31 127 -25 161
rect -71 89 -25 127
rect -71 55 -65 89
rect -31 55 -25 89
rect -71 17 -25 55
rect -71 -17 -65 17
rect -31 -17 -25 17
rect -71 -55 -25 -17
rect -71 -89 -65 -55
rect -31 -89 -25 -55
rect -71 -127 -25 -89
rect -71 -161 -65 -127
rect -31 -161 -25 -127
rect -71 -199 -25 -161
rect -71 -233 -65 -199
rect -31 -233 -25 -199
rect -71 -271 -25 -233
rect -71 -305 -65 -271
rect -31 -305 -25 -271
rect -71 -343 -25 -305
rect -71 -377 -65 -343
rect -31 -377 -25 -343
rect -71 -415 -25 -377
rect -71 -449 -65 -415
rect -31 -449 -25 -415
rect -71 -487 -25 -449
rect -71 -521 -65 -487
rect -31 -521 -25 -487
rect -71 -559 -25 -521
rect -71 -593 -65 -559
rect -31 -593 -25 -559
rect -71 -631 -25 -593
rect -71 -665 -65 -631
rect -31 -665 -25 -631
rect -71 -703 -25 -665
rect -71 -737 -65 -703
rect -31 -737 -25 -703
rect -71 -775 -25 -737
rect -71 -809 -65 -775
rect -31 -809 -25 -775
rect -71 -847 -25 -809
rect -71 -881 -65 -847
rect -31 -881 -25 -847
rect -71 -919 -25 -881
rect -71 -953 -65 -919
rect -31 -953 -25 -919
rect -71 -1000 -25 -953
rect 25 953 71 1000
rect 25 919 31 953
rect 65 919 71 953
rect 25 881 71 919
rect 25 847 31 881
rect 65 847 71 881
rect 25 809 71 847
rect 25 775 31 809
rect 65 775 71 809
rect 25 737 71 775
rect 25 703 31 737
rect 65 703 71 737
rect 25 665 71 703
rect 25 631 31 665
rect 65 631 71 665
rect 25 593 71 631
rect 25 559 31 593
rect 65 559 71 593
rect 25 521 71 559
rect 25 487 31 521
rect 65 487 71 521
rect 25 449 71 487
rect 25 415 31 449
rect 65 415 71 449
rect 25 377 71 415
rect 25 343 31 377
rect 65 343 71 377
rect 25 305 71 343
rect 25 271 31 305
rect 65 271 71 305
rect 25 233 71 271
rect 25 199 31 233
rect 65 199 71 233
rect 25 161 71 199
rect 25 127 31 161
rect 65 127 71 161
rect 25 89 71 127
rect 25 55 31 89
rect 65 55 71 89
rect 25 17 71 55
rect 25 -17 31 17
rect 65 -17 71 17
rect 25 -55 71 -17
rect 25 -89 31 -55
rect 65 -89 71 -55
rect 25 -127 71 -89
rect 25 -161 31 -127
rect 65 -161 71 -127
rect 25 -199 71 -161
rect 25 -233 31 -199
rect 65 -233 71 -199
rect 25 -271 71 -233
rect 25 -305 31 -271
rect 65 -305 71 -271
rect 25 -343 71 -305
rect 25 -377 31 -343
rect 65 -377 71 -343
rect 25 -415 71 -377
rect 25 -449 31 -415
rect 65 -449 71 -415
rect 25 -487 71 -449
rect 25 -521 31 -487
rect 65 -521 71 -487
rect 25 -559 71 -521
rect 25 -593 31 -559
rect 65 -593 71 -559
rect 25 -631 71 -593
rect 25 -665 31 -631
rect 65 -665 71 -631
rect 25 -703 71 -665
rect 25 -737 31 -703
rect 65 -737 71 -703
rect 25 -775 71 -737
rect 25 -809 31 -775
rect 65 -809 71 -775
rect 25 -847 71 -809
rect 25 -881 31 -847
rect 65 -881 71 -847
rect 25 -919 71 -881
rect 25 -953 31 -919
rect 65 -953 71 -919
rect 25 -1000 71 -953
rect 121 953 167 1000
rect 121 919 127 953
rect 161 919 167 953
rect 121 881 167 919
rect 121 847 127 881
rect 161 847 167 881
rect 121 809 167 847
rect 121 775 127 809
rect 161 775 167 809
rect 121 737 167 775
rect 121 703 127 737
rect 161 703 167 737
rect 121 665 167 703
rect 121 631 127 665
rect 161 631 167 665
rect 121 593 167 631
rect 121 559 127 593
rect 161 559 167 593
rect 121 521 167 559
rect 121 487 127 521
rect 161 487 167 521
rect 121 449 167 487
rect 121 415 127 449
rect 161 415 167 449
rect 121 377 167 415
rect 121 343 127 377
rect 161 343 167 377
rect 121 305 167 343
rect 121 271 127 305
rect 161 271 167 305
rect 121 233 167 271
rect 121 199 127 233
rect 161 199 167 233
rect 121 161 167 199
rect 121 127 127 161
rect 161 127 167 161
rect 121 89 167 127
rect 121 55 127 89
rect 161 55 167 89
rect 121 17 167 55
rect 121 -17 127 17
rect 161 -17 167 17
rect 121 -55 167 -17
rect 121 -89 127 -55
rect 161 -89 167 -55
rect 121 -127 167 -89
rect 121 -161 127 -127
rect 161 -161 167 -127
rect 121 -199 167 -161
rect 121 -233 127 -199
rect 161 -233 167 -199
rect 121 -271 167 -233
rect 121 -305 127 -271
rect 161 -305 167 -271
rect 121 -343 167 -305
rect 121 -377 127 -343
rect 161 -377 167 -343
rect 121 -415 167 -377
rect 121 -449 127 -415
rect 161 -449 167 -415
rect 121 -487 167 -449
rect 121 -521 127 -487
rect 161 -521 167 -487
rect 121 -559 167 -521
rect 121 -593 127 -559
rect 161 -593 167 -559
rect 121 -631 167 -593
rect 121 -665 127 -631
rect 161 -665 167 -631
rect 121 -703 167 -665
rect 121 -737 127 -703
rect 161 -737 167 -703
rect 121 -775 167 -737
rect 121 -809 127 -775
rect 161 -809 167 -775
rect 121 -847 167 -809
rect 121 -881 127 -847
rect 161 -881 167 -847
rect 121 -919 167 -881
rect 121 -953 127 -919
rect 161 -953 167 -919
rect 121 -1000 167 -953
<< end >>
