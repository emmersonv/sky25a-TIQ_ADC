magic
tech sky130A
magscale 1 2
timestamp 1755919380
<< nwell >>
rect -36 502 182 730
rect -16 478 152 502
rect 12 444 46 478
<< psubdiff >>
rect -80 -68 182 -28
rect -80 -104 -62 -68
rect -26 -104 30 -68
rect 66 -104 122 -68
rect 158 -104 182 -68
rect -80 -160 182 -104
rect -80 -196 -62 -160
rect -26 -196 30 -160
rect 66 -196 122 -160
rect 158 -196 182 -160
rect -80 -228 182 -196
<< nsubdiff >>
rect 0 664 146 694
rect 0 628 28 664
rect 64 628 146 664
rect 0 572 146 628
rect 0 536 28 572
rect 64 536 146 572
rect 0 494 146 536
<< psubdiffcont >>
rect -62 -104 -26 -68
rect 30 -104 66 -68
rect 122 -104 158 -68
rect -62 -196 -26 -160
rect 30 -196 66 -160
rect 122 -196 158 -160
<< nsubdiffcont >>
rect 28 628 64 664
rect 28 536 64 572
<< poly >>
rect -80 188 -14 204
rect 58 188 88 214
rect -80 152 -64 188
rect -30 152 88 188
rect -80 148 88 152
rect -80 136 -14 148
rect 58 136 88 148
<< polycont >>
rect -64 152 -30 188
<< locali >>
rect -80 664 182 680
rect -80 628 -64 664
rect -28 628 28 664
rect 64 628 120 664
rect 156 628 182 664
rect -80 572 182 628
rect -80 536 -64 572
rect -28 536 28 572
rect 64 536 120 572
rect 156 536 182 572
rect -80 508 182 536
rect 12 444 46 508
rect -80 188 -14 204
rect -80 152 -64 188
rect -30 152 -14 188
rect -80 136 -14 152
rect 100 188 134 236
rect 100 148 182 188
rect 100 114 134 148
rect 12 -44 46 22
rect -80 -68 182 -44
rect -80 -104 -62 -68
rect -26 -104 30 -68
rect 66 -104 122 -68
rect 158 -104 182 -68
rect -80 -160 182 -104
rect -80 -196 -62 -160
rect -26 -196 30 -160
rect 66 -196 122 -160
rect 158 -196 182 -160
rect -80 -212 182 -196
<< viali >>
rect -64 628 -28 664
rect 28 628 64 664
rect 120 628 156 664
rect -64 536 -28 572
rect 28 536 64 572
rect 120 536 156 572
rect -62 -104 -26 -68
rect 30 -104 66 -68
rect 122 -104 158 -68
rect -62 -196 -26 -160
rect 30 -196 66 -160
rect 122 -196 158 -160
<< metal1 >>
rect -80 664 182 680
rect -80 628 -64 664
rect -28 628 28 664
rect 64 628 120 664
rect 156 628 182 664
rect -80 572 182 628
rect -80 536 -64 572
rect -28 536 28 572
rect 64 536 120 572
rect 156 536 182 572
rect -80 508 182 536
rect -80 -68 182 -44
rect -80 -104 -62 -68
rect -26 -104 30 -68
rect 66 -104 122 -68
rect 158 -104 182 -68
rect -80 -160 182 -104
rect -80 -196 -62 -160
rect -26 -196 30 -160
rect 66 -196 122 -160
rect 158 -196 182 -160
rect -80 -212 182 -196
use sky130_fd_pr__nfet_01v8_PNPQML  sky130_fd_pr__nfet_01v8_PNPQML_0
timestamp 1755919380
transform 1 0 73 0 1 68
box -73 -68 73 68
use sky130_fd_pr__pfet_01v8_TH65V5  sky130_fd_pr__pfet_01v8_TH65V5_0
timestamp 1755919380
transform 1 0 73 0 1 340
box -109 -162 109 162
<< end >>
