magic
tech sky130A
magscale 1 2
timestamp 1756008383
<< error_s >>
rect -248 318 -232 470
rect -196 318 22 572
rect 212 318 430 572
rect 466 318 482 470
rect -232 302 22 318
rect 466 302 634 318
<< nwell >>
rect -196 2418 430 2646
rect -148 2410 -114 2418
rect 44 2410 78 2418
rect 156 2410 190 2418
rect 348 2410 382 2418
rect -196 2394 430 2410
rect -148 2360 -114 2394
rect 44 2360 78 2394
rect 156 2360 190 2394
rect 348 2360 382 2394
rect -248 302 -232 318
rect 28 300 206 330
rect 466 302 482 318
<< pwell >>
rect -274 -1376 496 -1124
<< psubdiff >>
rect -248 -1183 470 -1150
rect -248 -1217 -235 -1183
rect -201 -1217 -143 -1183
rect -109 -1217 -51 -1183
rect -17 -1217 41 -1183
rect 75 -1217 133 -1183
rect 167 -1217 225 -1183
rect 259 -1217 317 -1183
rect 351 -1217 409 -1183
rect 443 -1217 470 -1183
rect -248 -1275 470 -1217
rect -248 -1309 -235 -1275
rect -201 -1309 -143 -1275
rect -109 -1309 -51 -1275
rect -17 -1309 41 -1275
rect 75 -1309 133 -1275
rect 167 -1309 225 -1275
rect 259 -1309 317 -1275
rect 351 -1309 409 -1275
rect 443 -1309 470 -1275
rect -248 -1350 470 -1309
<< nsubdiff >>
rect -160 2579 394 2610
rect -160 2545 -109 2579
rect -75 2545 -17 2579
rect 17 2545 75 2579
rect 109 2545 167 2579
rect 201 2545 259 2579
rect 293 2545 351 2579
rect 385 2545 394 2579
rect -160 2487 394 2545
rect -160 2453 -109 2487
rect -75 2453 -17 2487
rect 17 2453 75 2487
rect 109 2453 167 2487
rect 201 2453 259 2487
rect 293 2453 351 2487
rect 385 2453 394 2487
rect -160 2410 394 2453
<< psubdiffcont >>
rect -235 -1217 -201 -1183
rect -143 -1217 -109 -1183
rect -51 -1217 -17 -1183
rect 41 -1217 75 -1183
rect 133 -1217 167 -1183
rect 225 -1217 259 -1183
rect 317 -1217 351 -1183
rect 409 -1217 443 -1183
rect -235 -1309 -201 -1275
rect -143 -1309 -109 -1275
rect -51 -1309 -17 -1275
rect 41 -1309 75 -1275
rect 133 -1309 167 -1275
rect 225 -1309 259 -1275
rect 317 -1309 351 -1275
rect 409 -1309 443 -1275
<< nsubdiffcont >>
rect -109 2545 -75 2579
rect -17 2545 17 2579
rect 75 2545 109 2579
rect 167 2545 201 2579
rect 259 2545 293 2579
rect 351 2545 385 2579
rect -109 2453 -75 2487
rect -17 2453 17 2487
rect 75 2453 109 2487
rect 167 2453 201 2487
rect 259 2453 293 2487
rect 351 2453 385 2487
<< poly >>
rect -248 326 -182 342
rect -248 292 -232 326
rect -198 306 -182 326
rect 28 306 206 330
rect -198 300 206 306
rect -198 292 332 300
rect -248 276 332 292
rect 58 252 88 276
<< polycont >>
rect -232 292 -198 326
<< locali >>
rect -248 2579 516 2596
rect -248 2545 -201 2579
rect -167 2545 -109 2579
rect -75 2545 -17 2579
rect 17 2545 75 2579
rect 109 2545 167 2579
rect 201 2545 259 2579
rect 293 2545 351 2579
rect 385 2545 516 2579
rect -248 2487 516 2545
rect -248 2453 -201 2487
rect -167 2453 -109 2487
rect -75 2453 -17 2487
rect 17 2453 75 2487
rect 109 2453 167 2487
rect 201 2453 259 2487
rect 293 2453 351 2487
rect 385 2453 516 2487
rect -248 2424 516 2453
rect -148 2360 -114 2424
rect 44 2360 78 2424
rect 156 2360 190 2424
rect 348 2360 382 2424
rect -248 326 -182 342
rect -248 292 -232 326
rect -198 292 -182 326
rect -248 276 -182 292
rect -52 316 -18 368
rect 252 316 286 352
rect 416 326 482 342
rect 416 316 432 326
rect -52 292 432 316
rect 466 292 482 326
rect -52 276 482 292
rect 100 230 134 276
rect 12 -1166 46 22
rect -248 -1183 470 -1166
rect -248 -1217 -235 -1183
rect -201 -1217 -143 -1183
rect -109 -1217 -51 -1183
rect -17 -1217 41 -1183
rect 75 -1217 133 -1183
rect 167 -1217 225 -1183
rect 259 -1217 317 -1183
rect 351 -1217 409 -1183
rect 443 -1217 470 -1183
rect -248 -1275 470 -1217
rect -248 -1309 -235 -1275
rect -201 -1309 -143 -1275
rect -109 -1309 -51 -1275
rect -17 -1309 41 -1275
rect 75 -1309 133 -1275
rect 167 -1309 225 -1275
rect 259 -1309 317 -1275
rect 351 -1309 409 -1275
rect 443 -1309 470 -1275
rect -248 -1334 470 -1309
<< viali >>
rect -201 2545 -167 2579
rect -109 2545 -75 2579
rect -17 2545 17 2579
rect 75 2545 109 2579
rect 167 2545 201 2579
rect 259 2545 293 2579
rect 351 2545 385 2579
rect -201 2453 -167 2487
rect -109 2453 -75 2487
rect -17 2453 17 2487
rect 75 2453 109 2487
rect 167 2453 201 2487
rect 259 2453 293 2487
rect 351 2453 385 2487
rect -232 292 -198 326
rect 432 292 466 326
rect -235 -1217 -201 -1183
rect -143 -1217 -109 -1183
rect -51 -1217 -17 -1183
rect 41 -1217 75 -1183
rect 133 -1217 167 -1183
rect 225 -1217 259 -1183
rect 317 -1217 351 -1183
rect 409 -1217 443 -1183
rect -235 -1309 -201 -1275
rect -143 -1309 -109 -1275
rect -51 -1309 -17 -1275
rect 41 -1309 75 -1275
rect 133 -1309 167 -1275
rect 225 -1309 259 -1275
rect 317 -1309 351 -1275
rect 409 -1309 443 -1275
<< metal1 >>
rect -248 2579 516 2596
rect -248 2545 -201 2579
rect -167 2545 -109 2579
rect -75 2545 -17 2579
rect 17 2545 75 2579
rect 109 2545 167 2579
rect 201 2545 259 2579
rect 293 2545 351 2579
rect 385 2545 516 2579
rect -248 2487 516 2545
rect -248 2453 -201 2487
rect -167 2453 -109 2487
rect -75 2453 -17 2487
rect 17 2453 75 2487
rect 109 2453 167 2487
rect 201 2453 259 2487
rect 293 2453 351 2487
rect 385 2453 516 2487
rect -248 2424 516 2453
rect -248 326 -182 342
rect -248 292 -232 326
rect -198 292 -182 326
rect -248 276 -182 292
rect 416 326 482 342
rect 416 292 432 326
rect 466 292 482 326
rect 416 276 482 292
rect -248 -1183 470 -1166
rect -248 -1217 -235 -1183
rect -201 -1217 -143 -1183
rect -109 -1217 -51 -1183
rect -17 -1217 41 -1183
rect 75 -1217 133 -1183
rect 167 -1217 225 -1183
rect 259 -1217 317 -1183
rect 351 -1217 409 -1183
rect 443 -1217 470 -1183
rect -248 -1275 470 -1217
rect -248 -1309 -235 -1275
rect -201 -1309 -143 -1275
rect -109 -1309 -51 -1275
rect -17 -1309 41 -1275
rect 75 -1309 133 -1275
rect 167 -1309 225 -1275
rect 259 -1309 317 -1275
rect 351 -1309 409 -1275
rect 443 -1309 470 -1275
rect -248 -1334 470 -1309
use sky130_fd_pr__nfet_01v8_QDUU3W  sky130_fd_pr__nfet_01v8_QDUU3W_0
timestamp 1756008383
transform 1 0 73 0 1 126
box -99 -126 99 126
use sky130_fd_pr__pfet_01v8_WELYR5  sky130_fd_pr__pfet_01v8_WELYR5_0
timestamp 1756008383
transform 1 0 -35 0 1 1356
box -161 -1062 161 1062
use sky130_fd_pr__pfet_01v8_WELYR5  sky130_fd_pr__pfet_01v8_WELYR5_1
timestamp 1756008383
transform 1 0 269 0 1 1356
box -161 -1062 161 1062
<< end >>
