magic
tech sky130A
magscale 1 2
timestamp 1756008383
<< nwell >>
rect -161 -862 161 862
<< pmos >>
rect -63 -800 -33 800
rect 33 -800 63 800
<< pdiff >>
rect -125 765 -63 800
rect -125 731 -113 765
rect -79 731 -63 765
rect -125 697 -63 731
rect -125 663 -113 697
rect -79 663 -63 697
rect -125 629 -63 663
rect -125 595 -113 629
rect -79 595 -63 629
rect -125 561 -63 595
rect -125 527 -113 561
rect -79 527 -63 561
rect -125 493 -63 527
rect -125 459 -113 493
rect -79 459 -63 493
rect -125 425 -63 459
rect -125 391 -113 425
rect -79 391 -63 425
rect -125 357 -63 391
rect -125 323 -113 357
rect -79 323 -63 357
rect -125 289 -63 323
rect -125 255 -113 289
rect -79 255 -63 289
rect -125 221 -63 255
rect -125 187 -113 221
rect -79 187 -63 221
rect -125 153 -63 187
rect -125 119 -113 153
rect -79 119 -63 153
rect -125 85 -63 119
rect -125 51 -113 85
rect -79 51 -63 85
rect -125 17 -63 51
rect -125 -17 -113 17
rect -79 -17 -63 17
rect -125 -51 -63 -17
rect -125 -85 -113 -51
rect -79 -85 -63 -51
rect -125 -119 -63 -85
rect -125 -153 -113 -119
rect -79 -153 -63 -119
rect -125 -187 -63 -153
rect -125 -221 -113 -187
rect -79 -221 -63 -187
rect -125 -255 -63 -221
rect -125 -289 -113 -255
rect -79 -289 -63 -255
rect -125 -323 -63 -289
rect -125 -357 -113 -323
rect -79 -357 -63 -323
rect -125 -391 -63 -357
rect -125 -425 -113 -391
rect -79 -425 -63 -391
rect -125 -459 -63 -425
rect -125 -493 -113 -459
rect -79 -493 -63 -459
rect -125 -527 -63 -493
rect -125 -561 -113 -527
rect -79 -561 -63 -527
rect -125 -595 -63 -561
rect -125 -629 -113 -595
rect -79 -629 -63 -595
rect -125 -663 -63 -629
rect -125 -697 -113 -663
rect -79 -697 -63 -663
rect -125 -731 -63 -697
rect -125 -765 -113 -731
rect -79 -765 -63 -731
rect -125 -800 -63 -765
rect -33 765 33 800
rect -33 731 -17 765
rect 17 731 33 765
rect -33 697 33 731
rect -33 663 -17 697
rect 17 663 33 697
rect -33 629 33 663
rect -33 595 -17 629
rect 17 595 33 629
rect -33 561 33 595
rect -33 527 -17 561
rect 17 527 33 561
rect -33 493 33 527
rect -33 459 -17 493
rect 17 459 33 493
rect -33 425 33 459
rect -33 391 -17 425
rect 17 391 33 425
rect -33 357 33 391
rect -33 323 -17 357
rect 17 323 33 357
rect -33 289 33 323
rect -33 255 -17 289
rect 17 255 33 289
rect -33 221 33 255
rect -33 187 -17 221
rect 17 187 33 221
rect -33 153 33 187
rect -33 119 -17 153
rect 17 119 33 153
rect -33 85 33 119
rect -33 51 -17 85
rect 17 51 33 85
rect -33 17 33 51
rect -33 -17 -17 17
rect 17 -17 33 17
rect -33 -51 33 -17
rect -33 -85 -17 -51
rect 17 -85 33 -51
rect -33 -119 33 -85
rect -33 -153 -17 -119
rect 17 -153 33 -119
rect -33 -187 33 -153
rect -33 -221 -17 -187
rect 17 -221 33 -187
rect -33 -255 33 -221
rect -33 -289 -17 -255
rect 17 -289 33 -255
rect -33 -323 33 -289
rect -33 -357 -17 -323
rect 17 -357 33 -323
rect -33 -391 33 -357
rect -33 -425 -17 -391
rect 17 -425 33 -391
rect -33 -459 33 -425
rect -33 -493 -17 -459
rect 17 -493 33 -459
rect -33 -527 33 -493
rect -33 -561 -17 -527
rect 17 -561 33 -527
rect -33 -595 33 -561
rect -33 -629 -17 -595
rect 17 -629 33 -595
rect -33 -663 33 -629
rect -33 -697 -17 -663
rect 17 -697 33 -663
rect -33 -731 33 -697
rect -33 -765 -17 -731
rect 17 -765 33 -731
rect -33 -800 33 -765
rect 63 765 125 800
rect 63 731 79 765
rect 113 731 125 765
rect 63 697 125 731
rect 63 663 79 697
rect 113 663 125 697
rect 63 629 125 663
rect 63 595 79 629
rect 113 595 125 629
rect 63 561 125 595
rect 63 527 79 561
rect 113 527 125 561
rect 63 493 125 527
rect 63 459 79 493
rect 113 459 125 493
rect 63 425 125 459
rect 63 391 79 425
rect 113 391 125 425
rect 63 357 125 391
rect 63 323 79 357
rect 113 323 125 357
rect 63 289 125 323
rect 63 255 79 289
rect 113 255 125 289
rect 63 221 125 255
rect 63 187 79 221
rect 113 187 125 221
rect 63 153 125 187
rect 63 119 79 153
rect 113 119 125 153
rect 63 85 125 119
rect 63 51 79 85
rect 113 51 125 85
rect 63 17 125 51
rect 63 -17 79 17
rect 113 -17 125 17
rect 63 -51 125 -17
rect 63 -85 79 -51
rect 113 -85 125 -51
rect 63 -119 125 -85
rect 63 -153 79 -119
rect 113 -153 125 -119
rect 63 -187 125 -153
rect 63 -221 79 -187
rect 113 -221 125 -187
rect 63 -255 125 -221
rect 63 -289 79 -255
rect 113 -289 125 -255
rect 63 -323 125 -289
rect 63 -357 79 -323
rect 113 -357 125 -323
rect 63 -391 125 -357
rect 63 -425 79 -391
rect 113 -425 125 -391
rect 63 -459 125 -425
rect 63 -493 79 -459
rect 113 -493 125 -459
rect 63 -527 125 -493
rect 63 -561 79 -527
rect 113 -561 125 -527
rect 63 -595 125 -561
rect 63 -629 79 -595
rect 113 -629 125 -595
rect 63 -663 125 -629
rect 63 -697 79 -663
rect 113 -697 125 -663
rect 63 -731 125 -697
rect 63 -765 79 -731
rect 113 -765 125 -731
rect 63 -800 125 -765
<< pdiffc >>
rect -113 731 -79 765
rect -113 663 -79 697
rect -113 595 -79 629
rect -113 527 -79 561
rect -113 459 -79 493
rect -113 391 -79 425
rect -113 323 -79 357
rect -113 255 -79 289
rect -113 187 -79 221
rect -113 119 -79 153
rect -113 51 -79 85
rect -113 -17 -79 17
rect -113 -85 -79 -51
rect -113 -153 -79 -119
rect -113 -221 -79 -187
rect -113 -289 -79 -255
rect -113 -357 -79 -323
rect -113 -425 -79 -391
rect -113 -493 -79 -459
rect -113 -561 -79 -527
rect -113 -629 -79 -595
rect -113 -697 -79 -663
rect -113 -765 -79 -731
rect -17 731 17 765
rect -17 663 17 697
rect -17 595 17 629
rect -17 527 17 561
rect -17 459 17 493
rect -17 391 17 425
rect -17 323 17 357
rect -17 255 17 289
rect -17 187 17 221
rect -17 119 17 153
rect -17 51 17 85
rect -17 -17 17 17
rect -17 -85 17 -51
rect -17 -153 17 -119
rect -17 -221 17 -187
rect -17 -289 17 -255
rect -17 -357 17 -323
rect -17 -425 17 -391
rect -17 -493 17 -459
rect -17 -561 17 -527
rect -17 -629 17 -595
rect -17 -697 17 -663
rect -17 -765 17 -731
rect 79 731 113 765
rect 79 663 113 697
rect 79 595 113 629
rect 79 527 113 561
rect 79 459 113 493
rect 79 391 113 425
rect 79 323 113 357
rect 79 255 113 289
rect 79 187 113 221
rect 79 119 113 153
rect 79 51 113 85
rect 79 -17 113 17
rect 79 -85 113 -51
rect 79 -153 113 -119
rect 79 -221 113 -187
rect 79 -289 113 -255
rect 79 -357 113 -323
rect 79 -425 113 -391
rect 79 -493 113 -459
rect 79 -561 113 -527
rect 79 -629 113 -595
rect 79 -697 113 -663
rect 79 -765 113 -731
<< poly >>
rect -63 800 -33 830
rect 33 800 63 830
rect -63 -826 -33 -800
rect 33 -826 63 -800
rect -63 -856 63 -826
<< locali >>
rect -113 773 -79 804
rect -113 701 -79 731
rect -113 629 -79 663
rect -113 561 -79 595
rect -113 493 -79 523
rect -113 425 -79 451
rect -113 357 -79 379
rect -113 289 -79 307
rect -113 221 -79 235
rect -113 153 -79 163
rect -113 85 -79 91
rect -113 17 -79 19
rect -113 -19 -79 -17
rect -113 -91 -79 -85
rect -113 -163 -79 -153
rect -113 -235 -79 -221
rect -113 -307 -79 -289
rect -113 -379 -79 -357
rect -113 -451 -79 -425
rect -113 -523 -79 -493
rect -113 -595 -79 -561
rect -113 -663 -79 -629
rect -113 -731 -79 -701
rect -113 -804 -79 -773
rect -17 773 17 804
rect -17 701 17 731
rect -17 629 17 663
rect -17 561 17 595
rect -17 493 17 523
rect -17 425 17 451
rect -17 357 17 379
rect -17 289 17 307
rect -17 221 17 235
rect -17 153 17 163
rect -17 85 17 91
rect -17 17 17 19
rect -17 -19 17 -17
rect -17 -91 17 -85
rect -17 -163 17 -153
rect -17 -235 17 -221
rect -17 -307 17 -289
rect -17 -379 17 -357
rect -17 -451 17 -425
rect -17 -523 17 -493
rect -17 -595 17 -561
rect -17 -663 17 -629
rect -17 -731 17 -701
rect -17 -804 17 -773
rect 79 773 113 804
rect 79 701 113 731
rect 79 629 113 663
rect 79 561 113 595
rect 79 493 113 523
rect 79 425 113 451
rect 79 357 113 379
rect 79 289 113 307
rect 79 221 113 235
rect 79 153 113 163
rect 79 85 113 91
rect 79 17 113 19
rect 79 -19 113 -17
rect 79 -91 113 -85
rect 79 -163 113 -153
rect 79 -235 113 -221
rect 79 -307 113 -289
rect 79 -379 113 -357
rect 79 -451 113 -425
rect 79 -523 113 -493
rect 79 -595 113 -561
rect 79 -663 113 -629
rect 79 -731 113 -701
rect 79 -804 113 -773
<< viali >>
rect -113 765 -79 773
rect -113 739 -79 765
rect -113 697 -79 701
rect -113 667 -79 697
rect -113 595 -79 629
rect -113 527 -79 557
rect -113 523 -79 527
rect -113 459 -79 485
rect -113 451 -79 459
rect -113 391 -79 413
rect -113 379 -79 391
rect -113 323 -79 341
rect -113 307 -79 323
rect -113 255 -79 269
rect -113 235 -79 255
rect -113 187 -79 197
rect -113 163 -79 187
rect -113 119 -79 125
rect -113 91 -79 119
rect -113 51 -79 53
rect -113 19 -79 51
rect -113 -51 -79 -19
rect -113 -53 -79 -51
rect -113 -119 -79 -91
rect -113 -125 -79 -119
rect -113 -187 -79 -163
rect -113 -197 -79 -187
rect -113 -255 -79 -235
rect -113 -269 -79 -255
rect -113 -323 -79 -307
rect -113 -341 -79 -323
rect -113 -391 -79 -379
rect -113 -413 -79 -391
rect -113 -459 -79 -451
rect -113 -485 -79 -459
rect -113 -527 -79 -523
rect -113 -557 -79 -527
rect -113 -629 -79 -595
rect -113 -697 -79 -667
rect -113 -701 -79 -697
rect -113 -765 -79 -739
rect -113 -773 -79 -765
rect -17 765 17 773
rect -17 739 17 765
rect -17 697 17 701
rect -17 667 17 697
rect -17 595 17 629
rect -17 527 17 557
rect -17 523 17 527
rect -17 459 17 485
rect -17 451 17 459
rect -17 391 17 413
rect -17 379 17 391
rect -17 323 17 341
rect -17 307 17 323
rect -17 255 17 269
rect -17 235 17 255
rect -17 187 17 197
rect -17 163 17 187
rect -17 119 17 125
rect -17 91 17 119
rect -17 51 17 53
rect -17 19 17 51
rect -17 -51 17 -19
rect -17 -53 17 -51
rect -17 -119 17 -91
rect -17 -125 17 -119
rect -17 -187 17 -163
rect -17 -197 17 -187
rect -17 -255 17 -235
rect -17 -269 17 -255
rect -17 -323 17 -307
rect -17 -341 17 -323
rect -17 -391 17 -379
rect -17 -413 17 -391
rect -17 -459 17 -451
rect -17 -485 17 -459
rect -17 -527 17 -523
rect -17 -557 17 -527
rect -17 -629 17 -595
rect -17 -697 17 -667
rect -17 -701 17 -697
rect -17 -765 17 -739
rect -17 -773 17 -765
rect 79 765 113 773
rect 79 739 113 765
rect 79 697 113 701
rect 79 667 113 697
rect 79 595 113 629
rect 79 527 113 557
rect 79 523 113 527
rect 79 459 113 485
rect 79 451 113 459
rect 79 391 113 413
rect 79 379 113 391
rect 79 323 113 341
rect 79 307 113 323
rect 79 255 113 269
rect 79 235 113 255
rect 79 187 113 197
rect 79 163 113 187
rect 79 119 113 125
rect 79 91 113 119
rect 79 51 113 53
rect 79 19 113 51
rect 79 -51 113 -19
rect 79 -53 113 -51
rect 79 -119 113 -91
rect 79 -125 113 -119
rect 79 -187 113 -163
rect 79 -197 113 -187
rect 79 -255 113 -235
rect 79 -269 113 -255
rect 79 -323 113 -307
rect 79 -341 113 -323
rect 79 -391 113 -379
rect 79 -413 113 -391
rect 79 -459 113 -451
rect 79 -485 113 -459
rect 79 -527 113 -523
rect 79 -557 113 -527
rect 79 -629 113 -595
rect 79 -697 113 -667
rect 79 -701 113 -697
rect 79 -765 113 -739
rect 79 -773 113 -765
<< metal1 >>
rect -119 773 -73 800
rect -119 739 -113 773
rect -79 739 -73 773
rect -119 701 -73 739
rect -119 667 -113 701
rect -79 667 -73 701
rect -119 629 -73 667
rect -119 595 -113 629
rect -79 595 -73 629
rect -119 557 -73 595
rect -119 523 -113 557
rect -79 523 -73 557
rect -119 485 -73 523
rect -119 451 -113 485
rect -79 451 -73 485
rect -119 413 -73 451
rect -119 379 -113 413
rect -79 379 -73 413
rect -119 341 -73 379
rect -119 307 -113 341
rect -79 307 -73 341
rect -119 269 -73 307
rect -119 235 -113 269
rect -79 235 -73 269
rect -119 197 -73 235
rect -119 163 -113 197
rect -79 163 -73 197
rect -119 125 -73 163
rect -119 91 -113 125
rect -79 91 -73 125
rect -119 53 -73 91
rect -119 19 -113 53
rect -79 19 -73 53
rect -119 -19 -73 19
rect -119 -53 -113 -19
rect -79 -53 -73 -19
rect -119 -91 -73 -53
rect -119 -125 -113 -91
rect -79 -125 -73 -91
rect -119 -163 -73 -125
rect -119 -197 -113 -163
rect -79 -197 -73 -163
rect -119 -235 -73 -197
rect -119 -269 -113 -235
rect -79 -269 -73 -235
rect -119 -307 -73 -269
rect -119 -341 -113 -307
rect -79 -341 -73 -307
rect -119 -379 -73 -341
rect -119 -413 -113 -379
rect -79 -413 -73 -379
rect -119 -451 -73 -413
rect -119 -485 -113 -451
rect -79 -485 -73 -451
rect -119 -523 -73 -485
rect -119 -557 -113 -523
rect -79 -557 -73 -523
rect -119 -595 -73 -557
rect -119 -629 -113 -595
rect -79 -629 -73 -595
rect -119 -667 -73 -629
rect -119 -701 -113 -667
rect -79 -701 -73 -667
rect -119 -739 -73 -701
rect -119 -773 -113 -739
rect -79 -773 -73 -739
rect -119 -800 -73 -773
rect -23 773 23 800
rect -23 739 -17 773
rect 17 739 23 773
rect -23 701 23 739
rect -23 667 -17 701
rect 17 667 23 701
rect -23 629 23 667
rect -23 595 -17 629
rect 17 595 23 629
rect -23 557 23 595
rect -23 523 -17 557
rect 17 523 23 557
rect -23 485 23 523
rect -23 451 -17 485
rect 17 451 23 485
rect -23 413 23 451
rect -23 379 -17 413
rect 17 379 23 413
rect -23 341 23 379
rect -23 307 -17 341
rect 17 307 23 341
rect -23 269 23 307
rect -23 235 -17 269
rect 17 235 23 269
rect -23 197 23 235
rect -23 163 -17 197
rect 17 163 23 197
rect -23 125 23 163
rect -23 91 -17 125
rect 17 91 23 125
rect -23 53 23 91
rect -23 19 -17 53
rect 17 19 23 53
rect -23 -19 23 19
rect -23 -53 -17 -19
rect 17 -53 23 -19
rect -23 -91 23 -53
rect -23 -125 -17 -91
rect 17 -125 23 -91
rect -23 -163 23 -125
rect -23 -197 -17 -163
rect 17 -197 23 -163
rect -23 -235 23 -197
rect -23 -269 -17 -235
rect 17 -269 23 -235
rect -23 -307 23 -269
rect -23 -341 -17 -307
rect 17 -341 23 -307
rect -23 -379 23 -341
rect -23 -413 -17 -379
rect 17 -413 23 -379
rect -23 -451 23 -413
rect -23 -485 -17 -451
rect 17 -485 23 -451
rect -23 -523 23 -485
rect -23 -557 -17 -523
rect 17 -557 23 -523
rect -23 -595 23 -557
rect -23 -629 -17 -595
rect 17 -629 23 -595
rect -23 -667 23 -629
rect -23 -701 -17 -667
rect 17 -701 23 -667
rect -23 -739 23 -701
rect -23 -773 -17 -739
rect 17 -773 23 -739
rect -23 -800 23 -773
rect 73 773 119 800
rect 73 739 79 773
rect 113 739 119 773
rect 73 701 119 739
rect 73 667 79 701
rect 113 667 119 701
rect 73 629 119 667
rect 73 595 79 629
rect 113 595 119 629
rect 73 557 119 595
rect 73 523 79 557
rect 113 523 119 557
rect 73 485 119 523
rect 73 451 79 485
rect 113 451 119 485
rect 73 413 119 451
rect 73 379 79 413
rect 113 379 119 413
rect 73 341 119 379
rect 73 307 79 341
rect 113 307 119 341
rect 73 269 119 307
rect 73 235 79 269
rect 113 235 119 269
rect 73 197 119 235
rect 73 163 79 197
rect 113 163 119 197
rect 73 125 119 163
rect 73 91 79 125
rect 113 91 119 125
rect 73 53 119 91
rect 73 19 79 53
rect 113 19 119 53
rect 73 -19 119 19
rect 73 -53 79 -19
rect 113 -53 119 -19
rect 73 -91 119 -53
rect 73 -125 79 -91
rect 113 -125 119 -91
rect 73 -163 119 -125
rect 73 -197 79 -163
rect 113 -197 119 -163
rect 73 -235 119 -197
rect 73 -269 79 -235
rect 113 -269 119 -235
rect 73 -307 119 -269
rect 73 -341 79 -307
rect 113 -341 119 -307
rect 73 -379 119 -341
rect 73 -413 79 -379
rect 113 -413 119 -379
rect 73 -451 119 -413
rect 73 -485 79 -451
rect 113 -485 119 -451
rect 73 -523 119 -485
rect 73 -557 79 -523
rect 113 -557 119 -523
rect 73 -595 119 -557
rect 73 -629 79 -595
rect 113 -629 119 -595
rect 73 -667 119 -629
rect 73 -701 79 -667
rect 113 -701 119 -667
rect 73 -739 119 -701
rect 73 -773 79 -739
rect 113 -773 119 -739
rect 73 -800 119 -773
<< end >>
