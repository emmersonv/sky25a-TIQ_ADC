magic
tech sky130A
magscale 1 2
timestamp 1756008383
<< nwell >>
rect -36 1490 894 3830
<< pwell >>
rect -62 -192 920 60
<< psubdiff >>
rect -36 1 894 34
rect -36 -33 31 1
rect 65 -33 123 1
rect 157 -33 215 1
rect 249 -33 307 1
rect 341 -33 399 1
rect 433 -33 491 1
rect 525 -33 583 1
rect 617 -33 675 1
rect 709 -33 767 1
rect 801 -33 894 1
rect -36 -91 894 -33
rect -36 -125 31 -91
rect 65 -125 123 -91
rect 157 -125 215 -91
rect 249 -125 307 -91
rect 341 -125 399 -91
rect 433 -125 491 -91
rect 525 -125 583 -91
rect 617 -125 675 -91
rect 709 -125 767 -91
rect 801 -125 894 -91
rect -36 -166 894 -125
<< nsubdiff >>
rect 0 3763 858 3794
rect 0 3729 65 3763
rect 99 3729 157 3763
rect 191 3729 249 3763
rect 283 3729 341 3763
rect 375 3729 433 3763
rect 467 3729 525 3763
rect 559 3729 617 3763
rect 651 3729 709 3763
rect 743 3729 801 3763
rect 835 3729 858 3763
rect 0 3671 858 3729
rect 0 3637 65 3671
rect 99 3637 157 3671
rect 191 3637 249 3671
rect 283 3637 341 3671
rect 375 3637 433 3671
rect 467 3637 525 3671
rect 559 3637 617 3671
rect 651 3637 709 3671
rect 743 3637 801 3671
rect 835 3637 858 3671
rect 0 3594 858 3637
<< psubdiffcont >>
rect 31 -33 65 1
rect 123 -33 157 1
rect 215 -33 249 1
rect 307 -33 341 1
rect 399 -33 433 1
rect 491 -33 525 1
rect 583 -33 617 1
rect 675 -33 709 1
rect 767 -33 801 1
rect 31 -125 65 -91
rect 123 -125 157 -91
rect 215 -125 249 -91
rect 307 -125 341 -91
rect 399 -125 433 -91
rect 491 -125 525 -91
rect 583 -125 617 -91
rect 675 -125 709 -91
rect 767 -125 801 -91
<< nsubdiffcont >>
rect 65 3729 99 3763
rect 157 3729 191 3763
rect 249 3729 283 3763
rect 341 3729 375 3763
rect 433 3729 467 3763
rect 525 3729 559 3763
rect 617 3729 651 3763
rect 709 3729 743 3763
rect 801 3729 835 3763
rect 65 3637 99 3671
rect 157 3637 191 3671
rect 249 3637 283 3671
rect 341 3637 375 3671
rect 433 3637 467 3671
rect 525 3637 559 3671
rect 617 3637 651 3671
rect 709 3637 743 3671
rect 801 3637 835 3671
<< poly >>
rect 0 1510 66 1526
rect 0 1476 16 1510
rect 50 1490 66 1510
rect 370 1490 400 1526
rect 50 1476 796 1490
rect 0 1460 796 1476
rect 188 1448 366 1460
rect 492 1448 670 1460
<< polycont >>
rect 16 1476 50 1510
<< locali >>
rect -36 3763 894 3780
rect -36 3729 65 3763
rect 99 3729 157 3763
rect 191 3729 249 3763
rect 283 3729 341 3763
rect 375 3729 433 3763
rect 467 3729 525 3763
rect 559 3729 617 3763
rect 651 3729 709 3763
rect 743 3729 801 3763
rect 835 3729 894 3763
rect -36 3671 894 3729
rect -36 3637 65 3671
rect 99 3637 157 3671
rect 191 3637 249 3671
rect 283 3637 341 3671
rect 375 3637 433 3671
rect 467 3637 525 3671
rect 559 3637 617 3671
rect 651 3637 709 3671
rect 743 3637 801 3671
rect 835 3637 894 3671
rect -36 3608 894 3637
rect 324 1650 358 3608
rect 0 1510 66 1526
rect 0 1476 16 1510
rect 50 1476 66 1510
rect 412 1500 446 1548
rect 792 1510 858 1526
rect 792 1500 808 1510
rect 0 1460 66 1476
rect 108 1476 808 1500
rect 842 1476 858 1510
rect 108 1460 858 1476
rect 108 1426 142 1460
rect 412 1426 446 1460
rect 716 1426 750 1460
rect 12 18 46 84
rect 204 18 238 84
rect 316 18 350 84
rect 508 18 542 84
rect 620 18 654 84
rect 812 18 846 84
rect -36 1 894 18
rect -36 -33 31 1
rect 65 -33 123 1
rect 157 -33 215 1
rect 249 -33 307 1
rect 341 -33 399 1
rect 433 -33 491 1
rect 525 -33 583 1
rect 617 -33 675 1
rect 709 -33 767 1
rect 801 -33 894 1
rect -36 -91 894 -33
rect -36 -125 31 -91
rect 65 -125 123 -91
rect 157 -125 215 -91
rect 249 -125 307 -91
rect 341 -125 399 -91
rect 433 -125 491 -91
rect 525 -125 583 -91
rect 617 -125 675 -91
rect 709 -125 767 -91
rect 801 -125 894 -91
rect -36 -150 894 -125
<< viali >>
rect 65 3729 99 3763
rect 157 3729 191 3763
rect 249 3729 283 3763
rect 341 3729 375 3763
rect 433 3729 467 3763
rect 525 3729 559 3763
rect 617 3729 651 3763
rect 709 3729 743 3763
rect 801 3729 835 3763
rect 65 3637 99 3671
rect 157 3637 191 3671
rect 249 3637 283 3671
rect 341 3637 375 3671
rect 433 3637 467 3671
rect 525 3637 559 3671
rect 617 3637 651 3671
rect 709 3637 743 3671
rect 801 3637 835 3671
rect 16 1476 50 1510
rect 808 1476 842 1510
rect 31 -33 65 1
rect 123 -33 157 1
rect 215 -33 249 1
rect 307 -33 341 1
rect 399 -33 433 1
rect 491 -33 525 1
rect 583 -33 617 1
rect 675 -33 709 1
rect 767 -33 801 1
rect 31 -125 65 -91
rect 123 -125 157 -91
rect 215 -125 249 -91
rect 307 -125 341 -91
rect 399 -125 433 -91
rect 491 -125 525 -91
rect 583 -125 617 -91
rect 675 -125 709 -91
rect 767 -125 801 -91
<< metal1 >>
rect -36 3763 894 3780
rect -36 3729 65 3763
rect 99 3729 157 3763
rect 191 3729 249 3763
rect 283 3729 341 3763
rect 375 3729 433 3763
rect 467 3729 525 3763
rect 559 3729 617 3763
rect 651 3729 709 3763
rect 743 3729 801 3763
rect 835 3729 894 3763
rect -36 3671 894 3729
rect -36 3637 65 3671
rect 99 3637 157 3671
rect 191 3637 249 3671
rect 283 3637 341 3671
rect 375 3637 433 3671
rect 467 3637 525 3671
rect 559 3637 617 3671
rect 651 3637 709 3671
rect 743 3637 801 3671
rect 835 3637 894 3671
rect -36 3608 894 3637
rect 0 1510 66 1526
rect 0 1476 16 1510
rect 50 1476 66 1510
rect 0 1460 66 1476
rect 792 1510 858 1526
rect 792 1476 808 1510
rect 842 1476 858 1510
rect 792 1460 858 1476
rect -36 1 894 18
rect -36 -33 31 1
rect 65 -33 123 1
rect 157 -33 215 1
rect 249 -33 307 1
rect 341 -33 399 1
rect 433 -33 491 1
rect 525 -33 583 1
rect 617 -33 675 1
rect 709 -33 767 1
rect 801 -33 894 1
rect -36 -91 894 -33
rect -36 -125 31 -91
rect 65 -125 123 -91
rect 157 -125 215 -91
rect 249 -125 307 -91
rect 341 -125 399 -91
rect 433 -125 491 -91
rect 525 -125 583 -91
rect 617 -125 675 -91
rect 709 -125 767 -91
rect 801 -125 894 -91
rect -36 -150 894 -125
use sky130_fd_pr__nfet_01v8_CTSNWR  sky130_fd_pr__nfet_01v8_CTSNWR_0
timestamp 1756008383
transform 1 0 125 0 1 755
box -151 -693 151 723
use sky130_fd_pr__nfet_01v8_CTSNWR  sky130_fd_pr__nfet_01v8_CTSNWR_1
timestamp 1756008383
transform 1 0 429 0 1 755
box -151 -693 151 723
use sky130_fd_pr__nfet_01v8_CTSNWR  sky130_fd_pr__nfet_01v8_CTSNWR_2
timestamp 1756008383
transform 1 0 733 0 1 755
box -151 -693 151 723
use sky130_fd_pr__pfet_01v8_FCTDLW  sky130_fd_pr__pfet_01v8_FCTDLW_0
timestamp 1756008383
transform 1 0 385 0 1 1599
box -109 -109 109 109
<< end >>
