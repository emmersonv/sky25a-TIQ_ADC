* NGSPICE file created from inverter_p0o5_n44.ext - technology: sky130A

.subckt sky130_fd_pr__nfet_01v8_3LP5BP a_63_n734# a_n33_n734# a_n63_n760# a_n125_n734#
+ VSUBS
X0 a_n33_n734# a_n63_n760# a_n125_n734# VSUBS sky130_fd_pr__nfet_01v8 ad=1.2111 pd=7.67 as=2.2754 ps=15.3 w=7.34 l=0.15
X1 a_63_n734# a_n63_n760# a_n33_n734# VSUBS sky130_fd_pr__nfet_01v8 ad=2.2754 pd=15.3 as=1.2111 ps=7.67 w=7.34 l=0.15
.ends

.subckt sky130_fd_pr__pfet_01v8_7SLTNL a_n15_n76# w_n109_n112# a_n73_n50# a_15_n50#
X0 a_15_n50# a_n15_n76# a_n73_n50# w_n109_n112# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.15
.ends

.subckt inverter_p0o5_n44 Vout Vin VDPWR VGND
Xsky130_fd_pr__nfet_01v8_3LP5BP_0 VGND Vout Vin VGND VGND sky130_fd_pr__nfet_01v8_3LP5BP
Xsky130_fd_pr__nfet_01v8_3LP5BP_1 VGND Vout Vin VGND VGND sky130_fd_pr__nfet_01v8_3LP5BP
Xsky130_fd_pr__nfet_01v8_3LP5BP_2 VGND Vout Vin VGND VGND sky130_fd_pr__nfet_01v8_3LP5BP
Xsky130_fd_pr__pfet_01v8_7SLTNL_0 Vin VDPWR VDPWR Vout sky130_fd_pr__pfet_01v8_7SLTNL
.ends

