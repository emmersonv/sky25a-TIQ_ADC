magic
tech sky130A
magscale 1 2
timestamp 1753650911
<< nmos >>
rect -63 -450 -33 450
rect 33 -450 63 450
<< ndiff >>
rect -125 438 -63 450
rect -125 -438 -113 438
rect -79 -438 -63 438
rect -125 -450 -63 -438
rect -33 438 33 450
rect -33 -438 -17 438
rect 17 -438 33 438
rect -33 -450 33 -438
rect 63 438 125 450
rect 63 -438 79 438
rect 113 -438 125 438
rect 63 -450 125 -438
<< ndiffc >>
rect -113 -438 -79 438
rect -17 -438 17 438
rect 79 -438 113 438
<< poly >>
rect -63 476 63 506
rect -63 450 -33 476
rect 33 450 63 476
rect -63 -476 -33 -450
rect 33 -476 63 -450
<< locali >>
rect -113 438 -79 454
rect -113 -454 -79 -438
rect -17 438 17 454
rect -17 -454 17 -438
rect 79 438 113 454
rect 79 -454 113 -438
<< viali >>
rect -113 -438 -79 438
rect -17 -438 17 438
rect 79 -438 113 438
<< metal1 >>
rect -119 438 -73 450
rect -119 -438 -113 438
rect -79 -438 -73 438
rect -119 -450 -73 -438
rect -23 438 23 450
rect -23 -438 -17 438
rect 17 -438 23 438
rect -23 -450 23 -438
rect 73 438 119 450
rect 73 -438 79 438
rect 113 -438 119 438
rect 73 -450 119 -438
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 4.5 l 0.150 m 1 nf 2 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 class mosfet compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
