magic
tech sky130A
magscale 1 2
timestamp 1755919380
<< error_s >>
rect 52 402 278 656
rect 166 394 278 402
rect 306 402 322 556
rect 306 388 474 402
<< nwell >>
rect -44 2116 278 2734
rect 4 2110 38 2116
rect 196 2110 230 2116
rect -44 2108 278 2110
rect 4 2060 38 2108
rect 196 2060 230 2108
rect 306 388 322 402
<< psubdiff >>
rect -88 -1094 322 -1062
rect -88 -1130 0 -1094
rect 36 -1130 92 -1094
rect 128 -1130 184 -1094
rect 220 -1130 276 -1094
rect 312 -1130 322 -1094
rect -88 -1186 322 -1130
rect -88 -1222 0 -1186
rect 36 -1222 92 -1186
rect 128 -1222 184 -1186
rect 220 -1222 276 -1186
rect 312 -1222 322 -1186
rect -88 -1262 322 -1222
<< nsubdiff >>
rect -8 2668 242 2698
rect -8 2632 34 2668
rect 70 2632 126 2668
rect 162 2632 242 2668
rect -8 2576 242 2632
rect -8 2540 34 2576
rect 70 2540 126 2576
rect 162 2540 242 2576
rect -8 2498 242 2540
<< psubdiffcont >>
rect 0 -1130 36 -1094
rect 92 -1130 128 -1094
rect 184 -1130 220 -1094
rect 276 -1130 312 -1094
rect 0 -1222 36 -1186
rect 92 -1222 128 -1186
rect 184 -1222 220 -1186
rect 276 -1222 312 -1186
<< nsubdiffcont >>
rect 34 2632 70 2668
rect 126 2632 162 2668
rect 34 2540 70 2576
rect 126 2540 162 2576
<< poly >>
rect -88 414 -22 430
rect -88 380 -72 414
rect -38 402 -22 414
rect -38 380 88 402
rect -88 364 88 380
rect 58 352 88 364
<< polycont >>
rect -72 380 -38 414
<< locali >>
rect -44 2668 278 2684
rect -44 2632 34 2668
rect 70 2632 126 2668
rect 162 2632 218 2668
rect 254 2632 278 2668
rect -44 2576 278 2632
rect -44 2540 34 2576
rect 70 2540 126 2576
rect 162 2540 218 2576
rect 254 2540 278 2576
rect -44 2512 278 2540
rect 4 2060 38 2512
rect 196 2060 230 2512
rect -88 414 -22 430
rect -88 380 -72 414
rect -38 380 -22 414
rect -88 364 -22 380
rect 100 404 134 452
rect 256 414 322 430
rect 256 404 272 414
rect 100 380 272 404
rect 306 380 322 414
rect 100 364 322 380
rect 100 330 134 364
rect 12 -1078 46 22
rect -88 -1094 322 -1078
rect -88 -1130 0 -1094
rect 36 -1130 92 -1094
rect 128 -1130 184 -1094
rect 220 -1130 276 -1094
rect 312 -1130 322 -1094
rect -88 -1186 322 -1130
rect -88 -1222 0 -1186
rect 36 -1222 92 -1186
rect 128 -1222 184 -1186
rect 220 -1222 276 -1186
rect 312 -1222 322 -1186
rect -88 -1246 322 -1222
<< viali >>
rect 34 2632 70 2668
rect 126 2632 162 2668
rect 218 2632 254 2668
rect 34 2540 70 2576
rect 126 2540 162 2576
rect 218 2540 254 2576
rect -72 380 -38 414
rect 272 380 306 414
rect 0 -1130 36 -1094
rect 92 -1130 128 -1094
rect 184 -1130 220 -1094
rect 276 -1130 312 -1094
rect 0 -1222 36 -1186
rect 92 -1222 128 -1186
rect 184 -1222 220 -1186
rect 276 -1222 312 -1186
<< metal1 >>
rect -44 2668 278 2684
rect -44 2632 34 2668
rect 70 2632 126 2668
rect 162 2632 218 2668
rect 254 2632 278 2668
rect -44 2576 278 2632
rect -44 2540 34 2576
rect 70 2540 126 2576
rect 162 2540 218 2576
rect 254 2540 278 2576
rect -44 2512 278 2540
rect -88 414 -22 430
rect -88 380 -72 414
rect -38 380 -22 414
rect -88 364 -22 380
rect 256 414 322 430
rect 256 380 272 414
rect 306 380 322 414
rect 256 364 322 380
rect -88 -1094 322 -1078
rect -88 -1130 0 -1094
rect 36 -1130 92 -1094
rect 128 -1130 184 -1094
rect 220 -1130 276 -1094
rect 312 -1130 322 -1094
rect -88 -1186 322 -1130
rect -88 -1222 0 -1186
rect 36 -1222 92 -1186
rect 128 -1222 184 -1186
rect 220 -1222 276 -1186
rect 312 -1222 322 -1186
rect -88 -1246 322 -1222
use sky130_fd_pr__nfet_01v8_PZUUQ8  sky130_fd_pr__nfet_01v8_PZUUQ8_0
timestamp 1755919380
transform 1 0 73 0 1 176
box -73 -176 73 176
use sky130_fd_pr__pfet_01v8_N885V5  sky130_fd_pr__pfet_01v8_N885V5_0
timestamp 1755919380
transform 1 0 117 0 1 1256
box -161 -862 161 862
<< end >>
