magic
tech sky130A
magscale 1 2
timestamp 1753144114
<< nwell >>
rect -36 1156 286 2308
<< psubdiff >>
rect -36 -14 286 34
rect -36 -118 34 -14
rect 216 -118 286 -14
rect -36 -166 286 -118
<< nsubdiff >>
rect 0 2224 250 2272
rect 0 2120 34 2224
rect 216 2120 250 2224
rect 0 2072 250 2120
<< psubdiffcont >>
rect 34 -118 216 -14
<< nsubdiffcont >>
rect 34 2120 216 2224
<< poly >>
rect -78 1176 -12 1192
rect -78 1142 -62 1176
rect -28 1156 -12 1176
rect 66 1156 96 1192
rect -28 1142 188 1156
rect -78 1126 188 1142
<< polycont >>
rect -62 1142 -28 1176
<< locali >>
rect 10 2224 240 2242
rect 10 2120 34 2224
rect 216 2120 240 2224
rect 10 2102 240 2120
rect 20 2022 54 2102
rect -78 1176 -12 1192
rect -78 1142 -62 1176
rect -28 1142 -12 1176
rect -78 1126 -12 1142
rect 108 1166 142 1214
rect 220 1176 286 1192
rect 220 1166 236 1176
rect 108 1142 236 1166
rect 270 1142 286 1176
rect 108 1126 286 1142
rect 108 1092 142 1126
rect 12 2 46 84
rect 204 2 238 84
rect 12 -14 238 2
rect 12 -118 34 -14
rect 216 -118 238 -14
rect 12 -134 238 -118
<< viali >>
rect 34 2120 216 2224
rect -62 1142 -28 1176
rect 236 1142 270 1176
rect 34 -118 216 -14
<< metal1 >>
rect 10 2224 240 2242
rect 10 2120 34 2224
rect 216 2120 240 2224
rect 10 2102 240 2120
rect -78 1176 -12 1192
rect -78 1142 -62 1176
rect -28 1142 -12 1176
rect -78 1126 -12 1142
rect 220 1176 286 1192
rect 220 1142 236 1176
rect 270 1142 286 1176
rect 220 1126 286 1142
rect 12 -14 238 2
rect 12 -118 34 -14
rect 216 -118 238 -14
rect 12 -134 238 -118
use sky130_fd_pr__nfet_01v8_QDUU3W  sky130_fd_pr__nfet_01v8_QDUU3W_0
timestamp 1753143363
transform 1 0 125 0 1 588
box -125 -526 125 556
use sky130_fd_pr__pfet_01v8_SDB5V5  sky130_fd_pr__pfet_01v8_SDB5V5_0
timestamp 1753143595
transform 1 0 81 0 1 1618
box -109 -462 109 462
<< labels >>
rlabel metal1 120 2224 136 2242 1 VDPWR
port 1 n
rlabel metal1 270 1156 286 1174 3 Vout
port 2 e
rlabel metal1 -78 1154 -62 1172 7 Vin
port 3 w
rlabel metal1 126 -134 140 -118 5 VGND
port 4 s
<< end >>
