magic
tech sky130A
magscale 1 2
timestamp 1756008383
<< error_s >>
rect 52 402 278 656
rect 306 402 322 556
rect 306 394 474 402
rect 322 388 474 394
<< nwell >>
rect -44 2116 278 2734
rect 4 2110 38 2116
rect 196 2110 230 2116
rect -44 2108 278 2110
rect 4 2060 38 2108
rect 196 2060 230 2108
rect 306 388 322 402
<< pwell >>
rect -114 -1288 348 -1036
<< psubdiff >>
rect -88 -1095 322 -1062
rect -88 -1129 1 -1095
rect 35 -1129 93 -1095
rect 127 -1129 185 -1095
rect 219 -1129 277 -1095
rect 311 -1129 322 -1095
rect -88 -1187 322 -1129
rect -88 -1221 1 -1187
rect 35 -1221 93 -1187
rect 127 -1221 185 -1187
rect 219 -1221 277 -1187
rect 311 -1221 322 -1187
rect -88 -1262 322 -1221
<< nsubdiff >>
rect -8 2667 242 2698
rect -8 2633 35 2667
rect 69 2633 127 2667
rect 161 2633 242 2667
rect -8 2575 242 2633
rect -8 2541 35 2575
rect 69 2541 127 2575
rect 161 2541 242 2575
rect -8 2498 242 2541
<< psubdiffcont >>
rect 1 -1129 35 -1095
rect 93 -1129 127 -1095
rect 185 -1129 219 -1095
rect 277 -1129 311 -1095
rect 1 -1221 35 -1187
rect 93 -1221 127 -1187
rect 185 -1221 219 -1187
rect 277 -1221 311 -1187
<< nsubdiffcont >>
rect 35 2633 69 2667
rect 127 2633 161 2667
rect 35 2541 69 2575
rect 127 2541 161 2575
<< poly >>
rect -88 414 -22 430
rect -88 380 -72 414
rect -38 402 -22 414
rect -38 380 88 402
rect -88 364 88 380
rect 58 352 88 364
<< polycont >>
rect -72 380 -38 414
<< locali >>
rect -44 2667 278 2684
rect -44 2633 35 2667
rect 69 2633 127 2667
rect 161 2633 219 2667
rect 253 2633 278 2667
rect -44 2575 278 2633
rect -44 2541 35 2575
rect 69 2541 127 2575
rect 161 2541 219 2575
rect 253 2541 278 2575
rect -44 2512 278 2541
rect 4 2060 38 2512
rect 196 2060 230 2512
rect -88 414 -22 430
rect -88 380 -72 414
rect -38 380 -22 414
rect -88 364 -22 380
rect 100 404 134 452
rect 256 414 322 430
rect 256 404 272 414
rect 100 380 272 404
rect 306 380 322 414
rect 100 364 322 380
rect 100 330 134 364
rect 12 -1078 46 22
rect -88 -1095 322 -1078
rect -88 -1129 1 -1095
rect 35 -1129 93 -1095
rect 127 -1129 185 -1095
rect 219 -1129 277 -1095
rect 311 -1129 322 -1095
rect -88 -1187 322 -1129
rect -88 -1221 1 -1187
rect 35 -1221 93 -1187
rect 127 -1221 185 -1187
rect 219 -1221 277 -1187
rect 311 -1221 322 -1187
rect -88 -1246 322 -1221
<< viali >>
rect 35 2633 69 2667
rect 127 2633 161 2667
rect 219 2633 253 2667
rect 35 2541 69 2575
rect 127 2541 161 2575
rect 219 2541 253 2575
rect -72 380 -38 414
rect 272 380 306 414
rect 1 -1129 35 -1095
rect 93 -1129 127 -1095
rect 185 -1129 219 -1095
rect 277 -1129 311 -1095
rect 1 -1221 35 -1187
rect 93 -1221 127 -1187
rect 185 -1221 219 -1187
rect 277 -1221 311 -1187
<< metal1 >>
rect -44 2667 278 2684
rect -44 2633 35 2667
rect 69 2633 127 2667
rect 161 2633 219 2667
rect 253 2633 278 2667
rect -44 2575 278 2633
rect -44 2541 35 2575
rect 69 2541 127 2575
rect 161 2541 219 2575
rect 253 2541 278 2575
rect -44 2512 278 2541
rect -88 414 -22 430
rect -88 380 -72 414
rect -38 380 -22 414
rect -88 364 -22 380
rect 256 414 322 430
rect 256 380 272 414
rect 306 380 322 414
rect 256 364 322 380
rect -88 -1095 322 -1078
rect -88 -1129 1 -1095
rect 35 -1129 93 -1095
rect 127 -1129 185 -1095
rect 219 -1129 277 -1095
rect 311 -1129 322 -1095
rect -88 -1187 322 -1129
rect -88 -1221 1 -1187
rect 35 -1221 93 -1187
rect 127 -1221 185 -1187
rect 219 -1221 277 -1187
rect 311 -1221 322 -1187
rect -88 -1246 322 -1221
use sky130_fd_pr__nfet_01v8_PZUUQ8  sky130_fd_pr__nfet_01v8_PZUUQ8_0
timestamp 1756008383
transform 1 0 73 0 1 176
box -99 -176 99 176
use sky130_fd_pr__pfet_01v8_N885V5  sky130_fd_pr__pfet_01v8_N885V5_0
timestamp 1756008383
transform 1 0 117 0 1 1256
box -161 -862 161 862
<< end >>
