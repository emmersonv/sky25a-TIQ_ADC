magic
tech sky130A
timestamp 1755919380
<< metal2 >>
rect 14151 1455 14168 3337
rect 14151 1438 14362 1455
rect 14324 280 14362 1438
rect 14324 252 14329 280
rect 14357 252 14362 280
rect 14324 247 14362 252
<< via2 >>
rect 14329 252 14357 280
<< metal3 >>
rect 8528 4188 8578 4197
rect 8528 4156 8537 4188
rect 8569 4156 8578 4188
rect 8528 992 8578 4156
rect 8712 4188 8762 4197
rect 8712 4156 8721 4188
rect 8753 4156 8762 4188
rect 8712 2216 8762 4156
rect 8962 4188 9012 4197
rect 8962 4156 8971 4188
rect 9003 4156 9012 4188
rect 8962 3440 9012 4156
rect 8712 2156 8963 2216
rect 8528 932 8962 992
rect 14322 280 15253 289
rect 14322 252 14329 280
rect 14357 252 15212 280
rect 14322 248 15212 252
rect 15244 248 15253 280
rect 14322 239 15253 248
<< via3 >>
rect 8537 4156 8569 4188
rect 8721 4156 8753 4188
rect 8971 4156 9003 4188
rect 15212 248 15244 280
<< metal4 >>
rect 3067 22476 3097 22576
rect 3343 22476 3373 22576
rect 3619 22476 3649 22576
rect 3895 22476 3925 22576
rect 4171 22476 4201 22576
rect 4447 22476 4477 22576
rect 4723 22476 4753 22576
rect 4999 22476 5029 22576
rect 5275 22476 5305 22576
rect 5551 22476 5581 22576
rect 5827 22476 5857 22576
rect 6103 22476 6133 22576
rect 6379 22476 6409 22576
rect 6655 22476 6685 22576
rect 6931 22476 6961 22576
rect 7207 22476 7237 22576
rect 7483 22476 7513 22576
rect 7759 22476 7789 22576
rect 8035 22476 8065 22576
rect 8311 22476 8341 22576
rect 8587 22476 8617 22576
rect 8863 22215 8893 22576
rect 8527 22185 8893 22215
rect 100 424 300 22076
rect 400 4077 600 22076
rect 8528 4188 8578 22185
rect 9139 22075 9169 22576
rect 8528 4156 8537 4188
rect 8569 4156 8578 4188
rect 8528 4147 8578 4156
rect 8712 22045 9169 22075
rect 8712 4188 8762 22045
rect 9415 21958 9445 22576
rect 9691 22476 9721 22576
rect 9967 22476 9997 22576
rect 10243 22476 10273 22576
rect 10519 22476 10549 22576
rect 10795 22476 10825 22576
rect 11071 22476 11101 22576
rect 11347 22476 11377 22576
rect 11623 22476 11653 22576
rect 11899 22476 11929 22576
rect 12175 22476 12205 22576
rect 12451 22476 12481 22576
rect 12727 22476 12757 22576
rect 13003 22476 13033 22576
rect 13279 22476 13309 22576
rect 13555 22476 13585 22576
rect 13831 22476 13861 22576
rect 14107 22476 14137 22576
rect 14383 22476 14413 22576
rect 14659 22476 14689 22576
rect 8712 4156 8721 4188
rect 8753 4156 8762 4188
rect 8712 4147 8762 4156
rect 8962 21928 9445 21958
rect 8962 4188 9012 21928
rect 8962 4156 8971 4188
rect 9003 4156 9012 4188
rect 8962 4147 9012 4156
rect 400 3875 11280 4077
rect 400 500 600 3875
rect 11120 3661 11280 3875
rect 10790 424 10950 632
rect 100 222 10950 424
rect 15181 280 15271 297
rect 15181 248 15212 280
rect 15244 248 15271 280
rect 1657 0 1747 100
rect 3589 0 3679 100
rect 5521 0 5611 100
rect 7453 0 7543 100
rect 9385 0 9475 100
rect 11317 0 11407 100
rect 13249 0 13339 100
rect 15181 0 15271 248
use full_tiq_adc_3  full_tiq_adc_3_0
timestamp 1755919380
transform 1 0 12720 0 1 422
box -3758 -38 2568 3432
<< labels >>
flabel metal4 s 14383 22476 14413 22576 0 FreeSans 300 90 0 0 clk
port 1 nsew
flabel metal4 s 14659 22476 14689 22576 0 FreeSans 300 90 0 0 ena
port 2 nsew
flabel metal4 s 14107 22476 14137 22576 0 FreeSans 300 90 0 0 rst_n
port 3 nsew
flabel metal4 s 15181 0 15271 100 0 FreeSans 600 0 0 0 ua[0]
port 4 nsew
flabel metal4 s 13249 0 13339 100 0 FreeSans 600 0 0 0 ua[1]
port 5 nsew
flabel metal4 s 11317 0 11407 100 0 FreeSans 600 0 0 0 ua[2]
port 6 nsew
flabel metal4 s 9385 0 9475 100 0 FreeSans 600 0 0 0 ua[3]
port 7 nsew
flabel metal4 s 7453 0 7543 100 0 FreeSans 600 0 0 0 ua[4]
port 8 nsew
flabel metal4 s 5521 0 5611 100 0 FreeSans 600 0 0 0 ua[5]
port 9 nsew
flabel metal4 s 3589 0 3679 100 0 FreeSans 600 0 0 0 ua[6]
port 10 nsew
flabel metal4 s 1657 0 1747 100 0 FreeSans 600 0 0 0 ua[7]
port 11 nsew
flabel metal4 s 13831 22476 13861 22576 0 FreeSans 300 90 0 0 ui_in[0]
port 12 nsew
flabel metal4 s 13555 22476 13585 22576 0 FreeSans 300 90 0 0 ui_in[1]
port 13 nsew
flabel metal4 s 13279 22476 13309 22576 0 FreeSans 300 90 0 0 ui_in[2]
port 14 nsew
flabel metal4 s 13003 22476 13033 22576 0 FreeSans 300 90 0 0 ui_in[3]
port 15 nsew
flabel metal4 s 12727 22476 12757 22576 0 FreeSans 300 90 0 0 ui_in[4]
port 16 nsew
flabel metal4 s 12451 22476 12481 22576 0 FreeSans 300 90 0 0 ui_in[5]
port 17 nsew
flabel metal4 s 12175 22476 12205 22576 0 FreeSans 300 90 0 0 ui_in[6]
port 18 nsew
flabel metal4 s 11899 22476 11929 22576 0 FreeSans 300 90 0 0 ui_in[7]
port 19 nsew
flabel metal4 s 11623 22476 11653 22576 0 FreeSans 300 90 0 0 uio_in[0]
port 20 nsew
flabel metal4 s 11347 22476 11377 22576 0 FreeSans 300 90 0 0 uio_in[1]
port 21 nsew
flabel metal4 s 11071 22476 11101 22576 0 FreeSans 300 90 0 0 uio_in[2]
port 22 nsew
flabel metal4 s 10795 22476 10825 22576 0 FreeSans 300 90 0 0 uio_in[3]
port 23 nsew
flabel metal4 s 10519 22476 10549 22576 0 FreeSans 300 90 0 0 uio_in[4]
port 24 nsew
flabel metal4 s 10243 22476 10273 22576 0 FreeSans 300 90 0 0 uio_in[5]
port 25 nsew
flabel metal4 s 9967 22476 9997 22576 0 FreeSans 300 90 0 0 uio_in[6]
port 26 nsew
flabel metal4 s 9691 22476 9721 22576 0 FreeSans 300 90 0 0 uio_in[7]
port 27 nsew
flabel metal4 s 4999 22476 5029 22576 0 FreeSans 300 90 0 0 uio_oe[0]
port 28 nsew
flabel metal4 s 4723 22476 4753 22576 0 FreeSans 300 90 0 0 uio_oe[1]
port 29 nsew
flabel metal4 s 4447 22476 4477 22576 0 FreeSans 300 90 0 0 uio_oe[2]
port 30 nsew
flabel metal4 s 4171 22476 4201 22576 0 FreeSans 300 90 0 0 uio_oe[3]
port 31 nsew
flabel metal4 s 3895 22476 3925 22576 0 FreeSans 300 90 0 0 uio_oe[4]
port 32 nsew
flabel metal4 s 3619 22476 3649 22576 0 FreeSans 300 90 0 0 uio_oe[5]
port 33 nsew
flabel metal4 s 3343 22476 3373 22576 0 FreeSans 300 90 0 0 uio_oe[6]
port 34 nsew
flabel metal4 s 3067 22476 3097 22576 0 FreeSans 300 90 0 0 uio_oe[7]
port 35 nsew
flabel metal4 s 7207 22476 7237 22576 0 FreeSans 300 90 0 0 uio_out[0]
port 36 nsew
flabel metal4 s 6931 22476 6961 22576 0 FreeSans 300 90 0 0 uio_out[1]
port 37 nsew
flabel metal4 s 6655 22476 6685 22576 0 FreeSans 300 90 0 0 uio_out[2]
port 38 nsew
flabel metal4 s 6379 22476 6409 22576 0 FreeSans 300 90 0 0 uio_out[3]
port 39 nsew
flabel metal4 s 6103 22476 6133 22576 0 FreeSans 300 90 0 0 uio_out[4]
port 40 nsew
flabel metal4 s 5827 22476 5857 22576 0 FreeSans 300 90 0 0 uio_out[5]
port 41 nsew
flabel metal4 s 5551 22476 5581 22576 0 FreeSans 300 90 0 0 uio_out[6]
port 42 nsew
flabel metal4 s 5275 22476 5305 22576 0 FreeSans 300 90 0 0 uio_out[7]
port 43 nsew
flabel metal4 s 9415 22476 9445 22576 0 FreeSans 300 90 0 0 uo_out[0]
port 44 nsew
flabel metal4 s 9139 22476 9169 22576 0 FreeSans 300 90 0 0 uo_out[1]
port 45 nsew
flabel metal4 s 8863 22476 8893 22576 0 FreeSans 300 90 0 0 uo_out[2]
port 46 nsew
flabel metal4 s 8587 22476 8617 22576 0 FreeSans 300 90 0 0 uo_out[3]
port 47 nsew
flabel metal4 s 8311 22476 8341 22576 0 FreeSans 300 90 0 0 uo_out[4]
port 48 nsew
flabel metal4 s 8035 22476 8065 22576 0 FreeSans 300 90 0 0 uo_out[5]
port 49 nsew
flabel metal4 s 7759 22476 7789 22576 0 FreeSans 300 90 0 0 uo_out[6]
port 50 nsew
flabel metal4 s 7483 22476 7513 22576 0 FreeSans 300 90 0 0 uo_out[7]
port 51 nsew
flabel metal4 s 100 500 300 22076 1 FreeSans 250 0 0 0 VDPWR
port 52 nsew
flabel metal4 s 400 500 600 22076 1 FreeSans 250 0 0 0 VGND
port 53 nsew
<< properties >>
string FIXED_BBOX 0 0 16100 22576
<< end >>
