* NGSPICE file created from inverter_p2_n18.ext - technology: sky130A

.subckt sky130_fd_pr__nfet_01v8_QQ9VTX a_63_n450# a_n63_n476# a_n33_n450# a_n125_n450#
+ VSUBS
X0 a_63_n450# a_n63_n476# a_n33_n450# VSUBS sky130_fd_pr__nfet_01v8 ad=1.395 pd=9.62 as=0.7425 ps=4.83 w=4.5 l=0.15
X1 a_n33_n450# a_n63_n476# a_n125_n450# VSUBS sky130_fd_pr__nfet_01v8 ad=0.7425 pd=4.83 as=1.395 ps=9.62 w=4.5 l=0.15
.ends

.subckt sky130_fd_pr__pfet_01v8_UCB5V5 a_15_n200# a_n15_n226# a_n73_n200# w_n109_n262#
X0 a_15_n200# a_n15_n226# a_n73_n200# w_n109_n262# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.15
.ends

.subckt inverter_p2_n18 VDPWR Vout Vin VGND
Xsky130_fd_pr__nfet_01v8_QQ9VTX_0 VGND Vin Vout VGND VGND sky130_fd_pr__nfet_01v8_QQ9VTX
Xsky130_fd_pr__nfet_01v8_QQ9VTX_1 VGND Vin Vout VGND VGND sky130_fd_pr__nfet_01v8_QQ9VTX
Xsky130_fd_pr__pfet_01v8_UCB5V5_0 Vout Vin VDPWR VDPWR sky130_fd_pr__pfet_01v8_UCB5V5
.ends

