magic
tech sky130A
magscale 1 2
timestamp 1756008383
<< error_s >>
rect -592 216 -576 366
rect -540 216 -322 470
rect -576 198 -322 216
<< nwell >>
rect -540 2312 678 2540
rect -512 2286 648 2312
rect -492 2254 -458 2286
rect -300 2254 -266 2286
rect 4 2254 38 2286
rect 196 2254 230 2286
rect 404 2254 438 2286
rect 596 2254 630 2286
rect -592 198 -576 216
<< pwell >>
rect -664 -1482 756 -1230
<< psubdiff >>
rect -638 -1289 730 -1256
rect -638 -1323 -607 -1289
rect -573 -1323 -515 -1289
rect -481 -1323 -423 -1289
rect -389 -1323 -331 -1289
rect -297 -1323 -239 -1289
rect -205 -1323 -147 -1289
rect -113 -1323 -55 -1289
rect -21 -1323 37 -1289
rect 71 -1323 129 -1289
rect 163 -1323 221 -1289
rect 255 -1323 313 -1289
rect 347 -1323 405 -1289
rect 439 -1323 497 -1289
rect 531 -1323 589 -1289
rect 623 -1323 681 -1289
rect 715 -1323 730 -1289
rect -638 -1381 730 -1323
rect -638 -1415 -607 -1381
rect -573 -1415 -515 -1381
rect -481 -1415 -423 -1381
rect -389 -1415 -331 -1381
rect -297 -1415 -239 -1381
rect -205 -1415 -147 -1381
rect -113 -1415 -55 -1381
rect -21 -1415 37 -1381
rect 71 -1415 129 -1381
rect 163 -1415 221 -1381
rect 255 -1415 313 -1381
rect 347 -1415 405 -1381
rect 439 -1415 497 -1381
rect 531 -1415 589 -1381
rect 623 -1415 681 -1381
rect 715 -1415 730 -1381
rect -638 -1456 730 -1415
<< nsubdiff >>
rect -504 2473 642 2504
rect -504 2439 -481 2473
rect -447 2439 -389 2473
rect -355 2439 -297 2473
rect -263 2439 -205 2473
rect -171 2439 -113 2473
rect -79 2439 -21 2473
rect 13 2439 71 2473
rect 105 2439 163 2473
rect 197 2439 255 2473
rect 289 2439 347 2473
rect 381 2439 439 2473
rect 473 2439 531 2473
rect 565 2439 642 2473
rect -504 2381 642 2439
rect -504 2347 -481 2381
rect -447 2347 -389 2381
rect -355 2347 -297 2381
rect -263 2347 -205 2381
rect -171 2347 -113 2381
rect -79 2347 -21 2381
rect 13 2347 71 2381
rect 105 2347 163 2381
rect 197 2347 255 2381
rect 289 2347 347 2381
rect 381 2347 439 2381
rect 473 2347 531 2381
rect 565 2347 642 2381
rect -504 2304 642 2347
<< psubdiffcont >>
rect -607 -1323 -573 -1289
rect -515 -1323 -481 -1289
rect -423 -1323 -389 -1289
rect -331 -1323 -297 -1289
rect -239 -1323 -205 -1289
rect -147 -1323 -113 -1289
rect -55 -1323 -21 -1289
rect 37 -1323 71 -1289
rect 129 -1323 163 -1289
rect 221 -1323 255 -1289
rect 313 -1323 347 -1289
rect 405 -1323 439 -1289
rect 497 -1323 531 -1289
rect 589 -1323 623 -1289
rect 681 -1323 715 -1289
rect -607 -1415 -573 -1381
rect -515 -1415 -481 -1381
rect -423 -1415 -389 -1381
rect -331 -1415 -297 -1381
rect -239 -1415 -205 -1381
rect -147 -1415 -113 -1381
rect -55 -1415 -21 -1381
rect 37 -1415 71 -1381
rect 129 -1415 163 -1381
rect 221 -1415 255 -1381
rect 313 -1415 347 -1381
rect 405 -1415 439 -1381
rect 497 -1415 531 -1381
rect 589 -1415 623 -1381
rect 681 -1415 715 -1381
<< nsubdiffcont >>
rect -481 2439 -447 2473
rect -389 2439 -355 2473
rect -297 2439 -263 2473
rect -205 2439 -171 2473
rect -113 2439 -79 2473
rect -21 2439 13 2473
rect 71 2439 105 2473
rect 163 2439 197 2473
rect 255 2439 289 2473
rect 347 2439 381 2473
rect 439 2439 473 2473
rect 531 2439 565 2473
rect -481 2347 -447 2381
rect -389 2347 -355 2381
rect -297 2347 -263 2381
rect -205 2347 -171 2381
rect -113 2347 -79 2381
rect -21 2347 13 2381
rect 71 2347 105 2381
rect 163 2347 197 2381
rect 255 2347 289 2381
rect 347 2347 381 2381
rect 439 2347 473 2381
rect 531 2347 565 2381
<< poly >>
rect -592 220 -526 236
rect -592 186 -576 220
rect -542 200 -526 220
rect -542 194 -394 200
rect -220 194 -42 224
rect 180 194 358 224
rect -542 186 580 194
rect -592 170 580 186
rect 58 146 88 170
<< polycont >>
rect -576 186 -542 220
<< locali >>
rect -592 2473 730 2490
rect -592 2439 -573 2473
rect -539 2439 -481 2473
rect -447 2439 -389 2473
rect -355 2439 -297 2473
rect -263 2439 -205 2473
rect -171 2439 -113 2473
rect -79 2439 -21 2473
rect 13 2439 71 2473
rect 105 2439 163 2473
rect 197 2439 255 2473
rect 289 2439 347 2473
rect 381 2439 439 2473
rect 473 2439 531 2473
rect 565 2439 623 2473
rect 657 2439 730 2473
rect -592 2381 730 2439
rect -592 2347 -573 2381
rect -539 2347 -481 2381
rect -447 2347 -389 2381
rect -355 2347 -297 2381
rect -263 2347 -205 2381
rect -171 2347 -113 2381
rect -79 2347 -21 2381
rect 13 2347 71 2381
rect 105 2347 163 2381
rect 197 2347 255 2381
rect 289 2347 347 2381
rect 381 2347 439 2381
rect 473 2347 531 2381
rect 565 2347 623 2381
rect 657 2347 730 2381
rect -592 2318 730 2347
rect -492 2254 -458 2318
rect -300 2254 -266 2318
rect 4 2254 38 2318
rect 196 2254 230 2318
rect 404 2254 438 2318
rect 596 2254 630 2318
rect -592 220 -526 236
rect -592 186 -576 220
rect -542 186 -526 220
rect -592 170 -526 186
rect -396 208 -362 246
rect -204 208 -170 246
rect -92 212 -58 246
rect 100 212 134 246
rect 308 212 342 246
rect 500 212 534 246
rect 664 222 730 238
rect 664 212 680 222
rect -92 208 680 212
rect -396 188 680 208
rect 714 188 730 222
rect -396 172 730 188
rect -396 170 -54 172
rect 100 124 134 172
rect 12 -1272 46 22
rect -638 -1289 730 -1272
rect -638 -1323 -607 -1289
rect -573 -1323 -515 -1289
rect -481 -1323 -423 -1289
rect -389 -1323 -331 -1289
rect -297 -1323 -239 -1289
rect -205 -1323 -147 -1289
rect -113 -1323 -55 -1289
rect -21 -1323 37 -1289
rect 71 -1323 129 -1289
rect 163 -1323 221 -1289
rect 255 -1323 313 -1289
rect 347 -1323 405 -1289
rect 439 -1323 497 -1289
rect 531 -1323 589 -1289
rect 623 -1323 681 -1289
rect 715 -1323 730 -1289
rect -638 -1381 730 -1323
rect -638 -1415 -607 -1381
rect -573 -1415 -515 -1381
rect -481 -1415 -423 -1381
rect -389 -1415 -331 -1381
rect -297 -1415 -239 -1381
rect -205 -1415 -147 -1381
rect -113 -1415 -55 -1381
rect -21 -1415 37 -1381
rect 71 -1415 129 -1381
rect 163 -1415 221 -1381
rect 255 -1415 313 -1381
rect 347 -1415 405 -1381
rect 439 -1415 497 -1381
rect 531 -1415 589 -1381
rect 623 -1415 681 -1381
rect 715 -1415 730 -1381
rect -638 -1440 730 -1415
<< viali >>
rect -573 2439 -539 2473
rect -481 2439 -447 2473
rect -389 2439 -355 2473
rect -297 2439 -263 2473
rect -205 2439 -171 2473
rect -113 2439 -79 2473
rect -21 2439 13 2473
rect 71 2439 105 2473
rect 163 2439 197 2473
rect 255 2439 289 2473
rect 347 2439 381 2473
rect 439 2439 473 2473
rect 531 2439 565 2473
rect 623 2439 657 2473
rect -573 2347 -539 2381
rect -481 2347 -447 2381
rect -389 2347 -355 2381
rect -297 2347 -263 2381
rect -205 2347 -171 2381
rect -113 2347 -79 2381
rect -21 2347 13 2381
rect 71 2347 105 2381
rect 163 2347 197 2381
rect 255 2347 289 2381
rect 347 2347 381 2381
rect 439 2347 473 2381
rect 531 2347 565 2381
rect 623 2347 657 2381
rect -576 186 -542 220
rect 680 188 714 222
rect -607 -1323 -573 -1289
rect -515 -1323 -481 -1289
rect -423 -1323 -389 -1289
rect -331 -1323 -297 -1289
rect -239 -1323 -205 -1289
rect -147 -1323 -113 -1289
rect -55 -1323 -21 -1289
rect 37 -1323 71 -1289
rect 129 -1323 163 -1289
rect 221 -1323 255 -1289
rect 313 -1323 347 -1289
rect 405 -1323 439 -1289
rect 497 -1323 531 -1289
rect 589 -1323 623 -1289
rect 681 -1323 715 -1289
rect -607 -1415 -573 -1381
rect -515 -1415 -481 -1381
rect -423 -1415 -389 -1381
rect -331 -1415 -297 -1381
rect -239 -1415 -205 -1381
rect -147 -1415 -113 -1381
rect -55 -1415 -21 -1381
rect 37 -1415 71 -1381
rect 129 -1415 163 -1381
rect 221 -1415 255 -1381
rect 313 -1415 347 -1381
rect 405 -1415 439 -1381
rect 497 -1415 531 -1381
rect 589 -1415 623 -1381
rect 681 -1415 715 -1381
<< metal1 >>
rect -592 2473 730 2490
rect -592 2439 -573 2473
rect -539 2439 -481 2473
rect -447 2439 -389 2473
rect -355 2439 -297 2473
rect -263 2439 -205 2473
rect -171 2439 -113 2473
rect -79 2439 -21 2473
rect 13 2439 71 2473
rect 105 2439 163 2473
rect 197 2439 255 2473
rect 289 2439 347 2473
rect 381 2439 439 2473
rect 473 2439 531 2473
rect 565 2439 623 2473
rect 657 2439 730 2473
rect -592 2381 730 2439
rect -592 2347 -573 2381
rect -539 2347 -481 2381
rect -447 2347 -389 2381
rect -355 2347 -297 2381
rect -263 2347 -205 2381
rect -171 2347 -113 2381
rect -79 2347 -21 2381
rect 13 2347 71 2381
rect 105 2347 163 2381
rect 197 2347 255 2381
rect 289 2347 347 2381
rect 381 2347 439 2381
rect 473 2347 531 2381
rect 565 2347 623 2381
rect 657 2347 730 2381
rect -592 2318 730 2347
rect -592 220 -526 236
rect -592 186 -576 220
rect -542 186 -526 220
rect -592 170 -526 186
rect 664 222 730 238
rect 664 188 680 222
rect 714 188 730 222
rect 664 172 730 188
rect -638 -1289 730 -1272
rect -638 -1323 -607 -1289
rect -573 -1323 -515 -1289
rect -481 -1323 -423 -1289
rect -389 -1323 -331 -1289
rect -297 -1323 -239 -1289
rect -205 -1323 -147 -1289
rect -113 -1323 -55 -1289
rect -21 -1323 37 -1289
rect 71 -1323 129 -1289
rect 163 -1323 221 -1289
rect 255 -1323 313 -1289
rect 347 -1323 405 -1289
rect 439 -1323 497 -1289
rect 531 -1323 589 -1289
rect 623 -1323 681 -1289
rect 715 -1323 730 -1289
rect -638 -1381 730 -1323
rect -638 -1415 -607 -1381
rect -573 -1415 -515 -1381
rect -481 -1415 -423 -1381
rect -389 -1415 -331 -1381
rect -297 -1415 -239 -1381
rect -205 -1415 -147 -1381
rect -113 -1415 -55 -1381
rect -21 -1415 37 -1381
rect 71 -1415 129 -1381
rect 163 -1415 221 -1381
rect 255 -1415 313 -1381
rect 347 -1415 405 -1381
rect 439 -1415 497 -1381
rect 531 -1415 589 -1381
rect 623 -1415 681 -1381
rect 715 -1415 730 -1381
rect -638 -1440 730 -1415
use sky130_fd_pr__nfet_01v8_PD6K7A  sky130_fd_pr__nfet_01v8_PD6K7A_0
timestamp 1756008383
transform 1 0 73 0 1 73
box -99 -73 99 73
use sky130_fd_pr__pfet_01v8_WGHLR5  sky130_fd_pr__pfet_01v8_WGHLR5_0
timestamp 1756008383
transform 1 0 -331 0 1 1250
box -209 -1062 209 1062
use sky130_fd_pr__pfet_01v8_WGHLR5  sky130_fd_pr__pfet_01v8_WGHLR5_1
timestamp 1756008383
transform 1 0 69 0 1 1250
box -209 -1062 209 1062
use sky130_fd_pr__pfet_01v8_WGHLR5  sky130_fd_pr__pfet_01v8_WGHLR5_2
timestamp 1756008383
transform 1 0 469 0 1 1250
box -209 -1062 209 1062
<< end >>
