magic
tech sky130A
magscale 1 2
timestamp 1753847028
<< nwell >>
rect -209 -1062 209 1062
<< pmos >>
rect -111 -1000 -81 1000
rect -15 -1000 15 1000
rect 81 -1000 111 1000
<< pdiff >>
rect -173 988 -111 1000
rect -173 -988 -161 988
rect -127 -988 -111 988
rect -173 -1000 -111 -988
rect -81 988 -15 1000
rect -81 -988 -65 988
rect -31 -988 -15 988
rect -81 -1000 -15 -988
rect 15 988 81 1000
rect 15 -988 31 988
rect 65 -988 81 988
rect 15 -1000 81 -988
rect 111 988 173 1000
rect 111 -988 127 988
rect 161 -988 173 988
rect 111 -1000 173 -988
<< pdiffc >>
rect -161 -988 -127 988
rect -65 -988 -31 988
rect 31 -988 65 988
rect 127 -988 161 988
<< poly >>
rect -111 1000 -81 1026
rect -15 1000 15 1026
rect 81 1000 111 1026
rect -111 -1026 -81 -1000
rect -15 -1026 15 -1000
rect 81 -1026 111 -1000
rect -111 -1056 111 -1026
<< locali >>
rect -161 988 -127 1004
rect -161 -1004 -127 -988
rect -65 988 -31 1004
rect -65 -1004 -31 -988
rect 31 988 65 1004
rect 31 -1004 65 -988
rect 127 988 161 1004
rect 127 -1004 161 -988
<< viali >>
rect -161 -988 -127 988
rect -65 -988 -31 988
rect 31 -988 65 988
rect 127 -988 161 988
<< metal1 >>
rect -167 988 -121 1000
rect -167 -988 -161 988
rect -127 -988 -121 988
rect -167 -1000 -121 -988
rect -71 988 -25 1000
rect -71 -988 -65 988
rect -31 -988 -25 988
rect -71 -1000 -25 -988
rect 25 988 71 1000
rect 25 -988 31 988
rect 65 -988 71 988
rect 25 -1000 71 -988
rect 121 988 167 1000
rect 121 -988 127 988
rect 161 -988 167 988
rect 121 -1000 167 -988
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 10 l 0.15 m 1 nf 3 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 class mosfet compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
