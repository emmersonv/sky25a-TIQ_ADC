magic
tech sky130A
magscale 1 2
timestamp 1755919380
<< error_s >>
rect 552 2760 554 2960
rect 588 2724 590 2996
<< nwell >>
rect -36 2172 588 2996
rect -36 656 590 2172
<< psubdiff >>
rect 0 -832 554 -800
rect 0 -868 20 -832
rect 56 -868 112 -832
rect 148 -868 204 -832
rect 240 -868 296 -832
rect 332 -868 388 -832
rect 424 -868 480 -832
rect 516 -868 554 -832
rect 0 -924 554 -868
rect 0 -960 20 -924
rect 56 -960 112 -924
rect 148 -960 204 -924
rect 240 -960 296 -924
rect 332 -960 388 -924
rect 424 -960 480 -924
rect 516 -960 554 -924
rect 0 -1000 554 -960
<< nsubdiff >>
rect 0 2930 554 2960
rect 0 2894 54 2930
rect 90 2894 146 2930
rect 182 2894 238 2930
rect 274 2894 330 2930
rect 366 2894 422 2930
rect 458 2894 554 2930
rect 0 2838 554 2894
rect 0 2802 54 2838
rect 90 2802 146 2838
rect 182 2802 238 2838
rect 274 2802 330 2838
rect 366 2802 422 2838
rect 458 2802 554 2838
rect 0 2760 554 2802
<< psubdiffcont >>
rect 20 -868 56 -832
rect 112 -868 148 -832
rect 204 -868 240 -832
rect 296 -868 332 -832
rect 388 -868 424 -832
rect 480 -868 516 -832
rect 20 -960 56 -924
rect 112 -960 148 -924
rect 204 -960 240 -924
rect 296 -960 332 -924
rect 388 -960 424 -924
rect 480 -960 516 -924
<< nsubdiffcont >>
rect 54 2894 90 2930
rect 146 2894 182 2930
rect 238 2894 274 2930
rect 330 2894 366 2930
rect 422 2894 458 2930
rect 54 2802 90 2838
rect 146 2802 182 2838
rect 238 2802 274 2838
rect 330 2802 366 2838
rect 422 2802 458 2838
<< poly >>
rect 0 676 66 692
rect 0 642 16 676
rect 50 656 66 676
rect 218 656 248 692
rect 50 644 492 656
rect 50 642 66 644
rect 0 626 66 642
rect 188 614 366 644
<< polycont >>
rect 16 642 50 676
<< locali >>
rect -36 2930 590 2946
rect -36 2894 54 2930
rect 90 2894 146 2930
rect 182 2894 238 2930
rect 274 2894 330 2930
rect 366 2894 422 2930
rect 458 2894 514 2930
rect 550 2894 590 2930
rect -36 2838 590 2894
rect -36 2802 54 2838
rect 90 2802 146 2838
rect 182 2802 238 2838
rect 274 2802 330 2838
rect 366 2802 422 2838
rect 458 2802 514 2838
rect 550 2802 590 2838
rect -36 2774 590 2802
rect 172 2106 206 2774
rect 0 676 66 692
rect 0 642 16 676
rect 50 642 66 676
rect 260 666 294 714
rect 488 676 554 692
rect 488 666 504 676
rect 0 626 66 642
rect 108 642 504 666
rect 538 642 554 676
rect 108 626 554 642
rect 108 576 142 626
rect 412 592 446 626
rect 12 -816 46 84
rect 204 -816 238 84
rect 316 -816 350 84
rect 508 -816 542 84
rect -36 -832 588 -816
rect -36 -868 20 -832
rect 56 -868 112 -832
rect 148 -868 204 -832
rect 240 -868 296 -832
rect 332 -868 388 -832
rect 424 -868 480 -832
rect 516 -868 588 -832
rect -36 -924 588 -868
rect -36 -960 20 -924
rect 56 -960 112 -924
rect 148 -960 204 -924
rect 240 -960 296 -924
rect 332 -960 388 -924
rect 424 -960 480 -924
rect 516 -960 588 -924
rect -36 -984 588 -960
<< viali >>
rect 54 2894 90 2930
rect 146 2894 182 2930
rect 238 2894 274 2930
rect 330 2894 366 2930
rect 422 2894 458 2930
rect 514 2894 550 2930
rect 54 2802 90 2838
rect 146 2802 182 2838
rect 238 2802 274 2838
rect 330 2802 366 2838
rect 422 2802 458 2838
rect 514 2802 550 2838
rect 16 642 50 676
rect 504 642 538 676
rect 20 -868 56 -832
rect 112 -868 148 -832
rect 204 -868 240 -832
rect 296 -868 332 -832
rect 388 -868 424 -832
rect 480 -868 516 -832
rect 20 -960 56 -924
rect 112 -960 148 -924
rect 204 -960 240 -924
rect 296 -960 332 -924
rect 388 -960 424 -924
rect 480 -960 516 -924
<< metal1 >>
rect -36 2930 590 2946
rect -36 2894 54 2930
rect 90 2894 146 2930
rect 182 2894 238 2930
rect 274 2894 330 2930
rect 366 2894 422 2930
rect 458 2894 514 2930
rect 550 2894 590 2930
rect -36 2838 590 2894
rect -36 2802 54 2838
rect 90 2802 146 2838
rect 182 2802 238 2838
rect 274 2802 330 2838
rect 366 2802 422 2838
rect 458 2802 514 2838
rect 550 2802 590 2838
rect -36 2774 590 2802
rect 0 676 66 692
rect 0 642 16 676
rect 50 642 66 676
rect 0 626 66 642
rect 488 676 554 692
rect 488 642 504 676
rect 538 642 554 676
rect 488 626 554 642
rect -36 -832 588 -816
rect -36 -868 20 -832
rect 56 -868 112 -832
rect 148 -868 204 -832
rect 240 -868 296 -832
rect 332 -868 388 -832
rect 424 -868 480 -832
rect 516 -868 588 -832
rect -36 -924 588 -868
rect -36 -960 20 -924
rect 56 -960 112 -924
rect 148 -960 204 -924
rect 240 -960 296 -924
rect 332 -960 388 -924
rect 424 -960 480 -924
rect 516 -960 588 -924
rect -36 -984 588 -960
use sky130_fd_pr__nfet_01v8_V2VUT3  sky130_fd_pr__nfet_01v8_V2VUT3_0
timestamp 1755919380
transform 1 0 125 0 1 338
box -125 -276 125 306
use sky130_fd_pr__nfet_01v8_V2VUT3  sky130_fd_pr__nfet_01v8_V2VUT3_1
timestamp 1755919380
transform 1 0 429 0 1 338
box -125 -276 125 306
use sky130_fd_pr__pfet_01v8_VGLYR5  sky130_fd_pr__pfet_01v8_VGLYR5_0
timestamp 1755919380
transform 1 0 233 0 1 1418
box -109 -762 109 762
<< end >>
