magic
tech sky130A
magscale 1 2
timestamp 1754087996
<< error_p >>
rect -161 -862 161 862
<< nwell >>
rect -161 -862 161 862
<< pmos >>
rect -63 -800 -33 800
rect 33 -800 63 800
<< pdiff >>
rect -125 788 -63 800
rect -125 -788 -113 788
rect -79 -788 -63 788
rect -125 -800 -63 -788
rect -33 788 33 800
rect -33 -788 -17 788
rect 17 -788 33 788
rect -33 -800 33 -788
rect 63 788 125 800
rect 63 -788 79 788
rect 113 -788 125 788
rect 63 -800 125 -788
<< pdiffc >>
rect -113 -788 -79 788
rect -17 -788 17 788
rect 79 -788 113 788
<< poly >>
rect -63 800 -33 830
rect 33 800 63 830
rect -63 -826 -33 -800
rect 33 -826 63 -800
rect -63 -856 63 -826
<< locali >>
rect -113 788 -79 804
rect -113 -804 -79 -788
rect -17 788 17 804
rect -17 -804 17 -788
rect 79 788 113 804
rect 79 -804 113 -788
<< viali >>
rect -113 -788 -79 788
rect -17 -788 17 788
rect 79 -788 113 788
<< metal1 >>
rect -119 788 -73 800
rect -119 -788 -113 788
rect -79 -788 -73 788
rect -119 -800 -73 -788
rect -23 788 23 800
rect -23 -788 -17 788
rect 17 -788 23 788
rect -23 -800 23 -788
rect 73 788 119 800
rect 73 -788 79 788
rect 113 -788 119 788
rect 73 -800 119 -788
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 8 l 0.15 m 1 nf 2 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 class mosfet compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
